* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
M_tn17 net3 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 SE net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net10 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 net5 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3_17 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tp17 net3 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net7 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net6 net3 net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net14 D net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 VDD SE net14 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp15 net1 cki net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp1_16 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS
