# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.97 1.79 6.08 1.79 6.08 2.12 3.97 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.98 1.83 3.655 1.83 3.655 2.35 6.355 2.35 6.355 1.79 7.25 1.79 7.25 2.195 6.615 2.195 6.615 2.68 3.395 2.68 3.395 2.09 2.98 2.09  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.939 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.785 2.75 1.785 2.75 2.12 0.28 2.12  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.45 3.095 2.45 3.095 3.05 6.845 3.05 6.845 2.445 7.5 2.445 7.5 1.56 3.77 1.56 3.77 0.99 4.11 0.99 4.11 1.22 6.01 1.22 6.01 0.99 6.35 0.99 6.35 1.22 7.7 1.22 7.73 1.22 7.73 2.675 7.7 2.675 7.075 2.675 7.075 3.28 2.865 3.28 2.865 2.68 1.595 2.68 1.595 3.335 1.365 3.335  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.995 0.575 2.995 0.575 3.62 2.385 3.62 2.385 2.995 2.615 2.995 2.615 3.62 7.305 3.62 7.305 2.995 7.535 2.995 7.535 3.62 7.7 3.62 8.4 3.62 8.4 4.22 7.7 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 1.595 0.3 1.595 1.015 1.365 1.015 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.635 0.475 0.635 0.475 1.31 2.485 1.31 2.485 0.53 7.7 0.53 7.7 0.76 2.715 0.76 2.715 1.545 0.245 1.545  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_2
