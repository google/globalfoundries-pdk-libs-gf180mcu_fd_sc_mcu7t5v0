* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_5 net_2 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 ZN C1 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_1 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_11 net_4 C2 VDD VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_10 VDD C1 net_4 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_8 net_4 B1 net_3 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_9 net_3 B2 net_4 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_7 ZN A2 net_3 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_6 net_3 A1 ZN VNW pfet_05v0 W=1.16e-06 L=5e-07
.ENDS
