# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 0.55 3.21 0.55 3.21 1.96 2.9 1.96  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 0.55 2.14 0.55 2.14 1.96 1.78 1.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.12 1.76 0.66 1.76 0.66 1.055 1.065 1.055 1.065 2.15 0.12 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3064 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 2.36 3.44 2.36 3.44 0.655 3.67 0.655 3.67 3.38 3.38 3.38 3.38 2.78 1.63 2.78 1.63 3.38 1.4 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.38 3.62 0.38 2.53 0.61 2.53 0.61 3.62 2.365 3.62 2.365 3.13 2.705 3.13 2.705 3.62 3.92 3.62 3.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.92 -0.3 3.92 0.3 0.61 0.3 0.61 0.805 0.38 0.805 0.38 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_1
