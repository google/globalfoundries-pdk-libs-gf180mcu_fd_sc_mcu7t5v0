* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_2_1 ZN A3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_1 VSS A4 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_0 ZN A4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0 VSS A3 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_1 VSS A1 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_0 ZN A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_6_1 net_2_1 A3 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD A4 net_2_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 net_2_0 A4 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 net_1_0 A3 net_2_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 net_0_1 A2 net_1_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 ZN A1 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 net_0_0 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 net_1 A2 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS
