# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.64 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.89 1.25 9.54 1.25 9.54 1.58 7.89 1.58  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 1.545 5.5 1.545 5.5 3.285 5.15 3.285  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.255 1.25 7.59 1.25 7.59 1.81 9.635 1.81 9.635 2.195 7.28 2.195 7.28 1.65 6.255 1.65  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 0.54 1.705 0.54 1.705 1.8 3.49 1.8 3.49 0.54 3.945 0.54 3.945 3.38 3.49 3.38 3.49 2.12 1.705 2.12 1.705 3.38 1.25 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.35 3.62 0.35 2.53 0.58 2.53 0.58 3.62 2.49 3.62 2.49 2.53 2.72 2.53 2.72 3.62 4.68 3.62 4.68 2.53 4.91 2.53 4.91 3.62 7.555 3.62 8.885 3.62 8.885 2.955 9.225 2.955 9.225 3.62 10.345 3.62 10.64 3.62 10.64 4.22 10.345 4.22 7.555 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.64 -0.3 10.64 0.3 9.17 0.3 9.17 0.835 8.94 0.835 8.94 0.3 5.01 0.3 5.01 0.835 4.78 0.835 4.78 0.3 2.77 0.3 2.77 0.835 2.54 0.835 2.54 0.3 0.53 0.3 0.53 0.835 0.3 0.835 0.3 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.985 2.965 7.555 2.965 7.555 3.195 5.755 3.195 5.755 1.315 4.47 1.315 4.47 1.78 4.24 1.78 4.24 1.085 5.755 1.085 5.755 0.55 7.115 0.55 7.115 0.78 5.985 0.78  ;
        POLYGON 6.615 1.96 6.955 1.96 6.955 2.49 10.005 2.49 10.005 0.54 10.345 0.54 10.345 3.39 9.96 3.39 9.96 2.725 6.615 2.725  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_4
