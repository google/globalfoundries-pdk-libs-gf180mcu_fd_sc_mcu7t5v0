# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.7 1.96 12.44 1.96 12.44 0.55 12.96 0.55 12.96 2.195 9.7 2.195  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.87 1.21 12.005 1.21 12.005 1.63 9.87 1.63  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.605 1.325 8.71 1.325 8.71 2.15 7.37 2.15 7.37 1.555 5.605 1.555  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.57 1.77 5.46 1.77 5.46 1.785 6.825 1.785 6.825 2.195 4.57 2.195  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.655 1.965 2.225 1.965 2.225 1.8 4.155 1.8 4.155 2.195 0.655 2.195  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.65 1.21 1.79 1.21 1.79 1.34 3.485 1.34 3.485 1.57 1.79 1.57 1.79 1.59 0.65 1.59  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.1688 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.225 0.74 2.25 0.74 2.25 0.865 4.925 0.865 4.925 0.845 5.265 0.845 5.265 0.865 9.05 0.865 9.05 0.79 9.47 0.79 9.47 2.44 13.255 2.44 13.255 0.57 13.485 0.57 13.485 2.67 9.05 2.67 9.05 1.095 2.02 1.095 2.02 0.97 0.225 0.97  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.225 3.62 0.225 2.53 0.565 2.53 0.565 3.62 2.32 3.62 2.32 3.04 2.55 3.04 2.55 3.62 4.36 3.62 4.36 3.04 4.59 3.04 4.59 3.62 13.55 3.62 14 3.62 14 4.22 13.55 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 14 -0.3 14 0.3 11.5 0.3 11.5 0.635 11.16 0.635 11.16 0.3 7.405 0.3 7.405 0.635 7.065 0.635 7.065 0.3 2.795 0.3 2.795 0.635 2.455 0.635 2.455 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.245 2.53 8.425 2.53 8.425 2.76 3.625 2.76 3.625 3.38 3.285 3.38 3.285 2.76 1.585 2.76 1.585 3.38 1.245 3.38  ;
        POLYGON 5.02 3.16 13.55 3.16 13.55 3.39 5.02 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_2
