# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.21 2.15 1.21 2.15 1.59 0.71 1.59  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.68 2.35 7.06 2.35 7.82 2.35 7.82 1.405 5.63 1.405 5.63 0.6 5.86 0.6 5.86 1.17 7.87 1.17 7.87 0.6 8.39 0.6 8.39 3.16 7.82 3.16 7.82 2.58 7.06 2.58 5.91 2.58 5.91 3.16 5.68 3.16  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.27 3.62 1.27 2.635 1.5 2.635 1.5 3.62 2.095 3.62 4.455 3.62 4.455 2.66 4.795 2.66 4.795 3.62 6.645 3.62 6.645 2.81 6.985 2.81 6.985 3.62 7.06 3.62 8.89 3.62 8.89 2.605 9.12 2.605 9.12 3.62 9.52 3.62 9.52 4.22 7.06 4.22 2.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.22 0.3 9.22 0.94 8.99 0.94 8.99 0.3 6.98 0.3 6.98 0.94 6.75 0.94 6.75 0.3 4.56 0.3 4.56 0.905 4.33 0.905 4.33 0.3 1.655 0.3 1.655 0.845 1.315 0.845 1.315 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 0.56 0.48 0.56 0.48 2.175 2.095 2.175 2.095 2.405 0.48 2.405 0.48 2.98 0.25 2.98  ;
        POLYGON 2.39 2.64 2.49 2.64 2.49 0.56 2.72 0.56 2.72 1.6 3.985 1.6 3.985 1.83 2.72 1.83 2.72 2.98 2.39 2.98  ;
        POLYGON 3.26 2.06 4.215 2.06 4.215 1.37 3.21 1.37 3.21 0.56 3.44 0.56 3.44 1.135 4.445 1.135 4.445 1.685 7.06 1.685 7.06 2.025 4.445 2.025 4.445 2.295 3.49 2.295 3.49 2.98 3.26 2.98  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_4
