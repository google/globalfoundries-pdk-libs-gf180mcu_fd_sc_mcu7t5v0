# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.08 1.55 9.31 1.55 9.31 1.79 12.05 1.79 12.05 2.12 9.08 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.57 1.225 12.05 1.225 12.05 1.56 9.57 1.56  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.125 1.91 5.65 1.91 5.65 1.8 7.815 1.8 7.815 2.14 4.125 2.14  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.525 1.785 3.04 1.785 3.04 1.45 5.39 1.45 5.39 1.68 3.27 1.68 3.27 2.15 0.525 2.15  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 1.325 2.58 1.325 2.58 0.99 6 0.99 6 1.21 8.31 1.21 8.31 1.56 5.77 1.56 5.77 1.22 2.81 1.22 2.81 1.555 0.87 1.555  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.496525 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.245 0.705 0.475 0.705 0.475 0.865 2.12 0.865 2.12 0.53 6.495 0.53 6.495 0.705 7.35 0.705 7.35 0.565 8.845 0.565 8.845 2.36 12.32 2.36 12.32 0.7 12.55 0.7 12.55 2.795 8.565 2.795 8.565 0.935 6.265 0.935 6.265 0.76 2.35 0.76 2.35 1.095 0.245 1.095  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.55 3.62 2.55 3.445 2.89 3.445 2.89 3.62 5.05 3.62 5.05 3.445 5.39 3.445 5.39 3.62 12.505 3.62 12.88 3.62 12.88 4.22 12.505 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 10.645 0.3 10.645 0.635 10.305 0.635 10.305 0.3 7.065 0.3 7.065 0.475 6.725 0.475 6.725 0.3 1.87 0.3 1.87 0.635 1.53 0.635 1.53 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.31 2.525 7.41 2.525 7.41 2.755 1.31 2.755  ;
        POLYGON 0.345 2.46 0.575 2.46 0.575 3.12 2.075 3.12 2.075 2.985 6.195 2.985 6.195 3.135 8.105 3.135 8.105 2.46 8.335 2.46 8.335 3.135 12.505 3.135 12.505 3.365 5.855 3.365 5.855 3.215 2.29 3.215 2.29 3.35 0.345 3.35  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_2
