# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.215 1.77 2.34 1.77 2.34 1.445 3.87 1.445 3.87 1.675 2.57 1.675 2.57 2.135 1.215 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.825 1.905 5.42 1.905 5.42 1.8 7.545 1.8 7.545 2.135 2.825 2.135  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.68 3.89 0.68 3.89 0.985 4.235 0.985 4.235 0.99 7.17 0.99 7.17 1.38 6.83 1.38 6.83 1.22 4.005 1.22 4.005 1.215 2.05 1.215 2.05 1.385 0.96 1.385  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.77 0.985 1.77 0.985 2.365 7.96 2.365 7.96 1.645 8.28 1.645 8.28 2.595 0.14 2.595  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.54 2.38 11.55 2.38 11.85 2.38 11.85 1.1 9.485 1.1 9.485 0.53 9.825 0.53 9.825 0.87 11.725 0.87 11.725 0.53 12.23 0.53 12.23 2.725 11.945 2.725 11.945 3.195 11.58 3.195 11.58 2.725 11.55 2.725 9.905 2.725 9.905 3.195 9.54 3.195  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.26 3.62 0.26 3.005 0.49 3.005 0.49 3.62 2.245 3.62 2.245 3.285 2.585 3.285 2.585 3.62 4.285 3.62 4.285 3.285 4.625 3.285 4.625 3.62 6.325 3.62 6.325 3.285 6.665 3.285 6.665 3.62 8.365 3.62 8.365 3.285 8.705 3.285 8.705 3.62 10.585 3.62 10.585 3.215 10.925 3.215 10.925 3.62 11.55 3.62 12.68 3.62 12.68 2.69 12.91 2.69 12.91 3.62 13.44 3.62 13.44 4.22 11.55 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 13.13 0.3 13.13 0.905 12.9 0.905 12.9 0.3 10.945 0.3 10.945 0.64 10.605 0.64 10.605 0.3 8.65 0.3 8.65 0.695 8.42 0.695 8.42 0.3 0.49 0.3 0.49 0.765 0.26 0.765 0.26 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.185 2.825 8.86 2.825 8.86 1.155 7.96 1.155 7.96 0.76 4.285 0.76 4.285 0.53 8.19 0.53 8.19 0.925 9.09 0.925 9.09 1.525 11.55 1.525 11.55 1.755 9.09 1.755 9.09 3.055 1.185 3.055  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_4
