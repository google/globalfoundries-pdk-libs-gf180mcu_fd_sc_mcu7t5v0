# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.965 1.79 3.27 1.79 3.27 2.12 0.965 2.12  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.78 1.24 4.045 1.24 4.045 2.795 3.5 2.795 3.5 1.56 0.78 1.56  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.38 1.8 7.38 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.64 2.11 10.935 2.11 11.3 2.11 11.3 1.38 10.64 1.38 10.64 0.555 11.1 0.555 11.1 1.13 11.66 1.13 11.66 2.34 11.1 2.34 11.1 3.38 10.935 3.38 10.64 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3 1.595 3 1.595 3.62 3.16 3.62 5.365 3.62 5.365 3 5.595 3 5.595 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 9.525 3.62 9.525 2.57 9.755 2.57 9.755 3.62 10.935 3.62 11.665 3.62 11.665 2.57 11.895 2.57 11.895 3.62 12.32 3.62 12.32 4.22 10.935 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.995 0.3 11.995 0.895 11.765 0.895 11.765 0.3 9.755 0.3 9.755 0.895 9.525 0.895 9.525 0.3 5.695 0.3 5.695 0.86 5.465 0.86 5.465 0.3 1.595 0.3 1.595 0.86 1.365 0.86 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 2.35 3.16 2.35 3.16 2.58 0.575 2.58 0.575 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 0.76 3.41 0.76 3.41 0.53 4.56 0.53 4.56 1.225 6.53 1.225 6.53 1.455 4.56 1.455 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.63 9.245 1.63 9.245 1.86 7.97 1.86 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 8.505 2.11 9.585 2.11 9.585 1.38 8.405 1.38 8.405 0.555 8.635 0.555 8.635 1.15 9.815 1.15 9.815 1.63 10.935 1.63 10.935 1.86 9.815 1.86 9.815 2.34 8.735 2.34 8.735 3.38 8.505 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_2
