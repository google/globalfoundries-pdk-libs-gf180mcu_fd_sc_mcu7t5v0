# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.54 1.77 1.25 1.77 1.25 1.12 1.57 1.12 1.57 2.15 0.54 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.8 1.12 2.12 1.12 2.12 2.415 1.8 2.415  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.36 1.12 2.91 1.12 2.91 2.415 2.36 2.415  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8756 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.57 0.65 5.01 0.65 5.01 3.38 4.57 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 3.285 1.55 3.285 1.55 3.62 3.745 3.62 3.745 2.53 3.975 2.53 3.975 3.62 4.315 3.62 5.6 3.62 5.6 4.22 4.315 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 3.875 0.3 3.875 1.09 3.645 1.09 3.645 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 2.825 3.185 2.825 3.185 0.805 0.53 0.805 0.53 1.035 0.19 1.035 0.19 0.575 3.415 0.575 3.415 1.46 4.315 1.46 4.315 1.8 3.415 1.8 3.415 3.055 2.57 3.055 2.57 3.34 2.23 3.34 2.23 3.055 0.53 3.055 0.53 3.34 0.19 3.34  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_1
