# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.37 1.74 1.95 1.74 1.95 2.15 0.37 2.15  ;
        POLYGON 3.035 1.74 4.315 1.74 4.315 2.15 3.035 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6096 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.71 2.39 3.835 2.39 3.835 3.39 3.605 3.39 3.605 2.77 1.595 2.77 1.595 3.39 1.365 3.39 1.365 2.39 2.33 2.39 2.33 1.44 1.365 1.44 1.365 0.675 1.595 0.675 1.595 1.06 3.605 1.06 3.605 0.675 3.835 0.675 3.835 1.44 2.71 1.44  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.615 0.475 2.615 0.475 3.62 2.485 3.62 2.485 3.13 2.715 3.13 2.715 3.62 4.725 3.62 4.725 2.62 4.955 2.62 4.955 3.62 5.6 3.62 5.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 0.975 4.725 0.975 4.725 0.3 2.715 0.3 2.715 0.775 2.485 0.775 2.485 0.3 0.475 0.3 0.475 0.97 0.245 0.97 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_4
