# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.1 1.685 1.33 1.685 1.33 2.015 3.905 2.015 3.905 1.8 5.845 1.8 5.845 2.015 10.47 2.015 10.47 2.245 1.1 2.245  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 1.2 3.965 1.2 3.965 1.305 6.585 1.305 6.585 1.555 7.62 1.555 7.62 1.785 6.355 1.785 6.355 1.57 3.47 1.57 3.47 1.775 1.64 1.775  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2701 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.17 1.035 13.56 1.035 13.56 1.77 15.9 1.77 15.9 1.035 16.24 1.035 16.24 2.885 15.85 2.885 15.85 2.15 13.51 2.15 13.51 2.885 13.17 2.885  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0903 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.22 2.245 19.86 2.245 20.25 2.245 20.25 1.37 18.22 1.37 18.22 0.54 18.605 0.54 18.605 1.135 20.25 1.135 20.25 0.65 20.845 0.65 20.845 3.39 20.25 3.39 20.25 2.48 19.86 2.48 18.56 2.48 18.56 3.39 18.22 3.39  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.145 0.475 3.145 0.475 3.62 2.335 3.62 2.335 3.105 2.565 3.105 2.565 3.62 4.425 3.62 4.425 3.105 4.655 3.105 4.655 3.62 8.3 3.62 8.3 3.445 8.64 3.445 8.64 3.62 12.045 3.62 12.045 3.285 12.385 3.285 12.385 3.62 14.51 3.62 14.51 3.285 14.85 3.285 14.85 3.62 17.125 3.62 17.125 2.73 17.355 2.73 17.355 3.62 19.395 3.62 19.395 2.73 19.625 2.73 19.625 3.62 19.86 3.62 21.605 3.62 21.605 2.73 21.835 2.73 21.835 3.62 22.4 3.62 22.4 4.22 19.86 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 21.965 0.3 21.965 0.935 21.735 0.935 21.735 0.3 19.78 0.3 19.78 0.735 19.44 0.735 19.44 0.3 17.455 0.3 17.455 0.935 17.225 0.935 17.225 0.3 14.9 0.3 14.9 0.635 14.56 0.635 14.56 0.3 12.44 0.3 12.44 1.12 12.09 1.12 12.09 0.3 4.71 0.3 4.71 1.075 4.37 1.075 4.37 0.3 0.475 0.3 0.475 0.69 0.245 0.69 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.72 0.63 11.1 0.63 11.1 1.075 10.76 1.075 10.76 0.86 8.64 0.86 8.64 0.915 8.3 0.915 8.3 0.86 6.06 0.86 6.06 1.075 5.72 1.075  ;
        POLYGON 0.87 2.525 10.7 2.525 10.7 1.815 12.88 1.815 12.88 2.045 10.93 2.045 10.93 2.755 3.69 2.755 3.69 3.39 3.35 3.39 3.35 2.815 1.6 2.815 1.6 3.39 1.255 3.39 1.255 2.815 0.64 2.815 0.64 1.09 1.025 1.09 1.025 0.54 2.67 0.54 2.67 0.77 1.255 0.77 1.255 1.32 0.87 1.32  ;
        POLYGON 5.72 2.985 11.385 2.985 11.385 2.825 12.89 2.825 12.89 3.115 13.825 3.115 13.825 2.75 15.545 2.75 15.545 3.115 16.47 3.115 16.47 0.76 15.565 0.76 15.565 1.235 14.03 1.235 14.03 0.76 12.92 0.76 12.92 1.585 9.64 1.585 9.64 1.38 7.885 1.38 7.885 1.325 6.84 1.325 6.84 1.09 8.115 1.09 8.115 1.145 9.64 1.145 9.64 1.09 9.98 1.09 9.98 1.35 12.69 1.35 12.69 0.53 14.26 0.53 14.26 1.005 15.335 1.005 15.335 0.53 16.7 0.53 16.7 1.74 19.86 1.74 19.86 1.97 16.7 1.97 16.7 3.345 15.315 3.345 15.315 2.98 14.055 2.98 14.055 3.345 12.66 3.345 12.66 3.055 11.615 3.055 11.615 3.215 5.72 3.215  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_4
