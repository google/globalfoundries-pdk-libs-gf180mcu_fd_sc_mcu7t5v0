* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyc_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_8 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_8 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_8 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2_36 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_8 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_8 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_8 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_16 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_32 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_16_16 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS
