# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.49 1.79 19.73 1.79 19.73 2.35 22.8 2.35 22.8 1.95 23.14 1.95 23.14 2.35 23.82 2.35 23.82 1.95 24.16 1.95 24.16 2.35 27.42 2.35 27.42 1.72 27.715 1.72 27.715 2.58 24.8 2.58 24.8 2.68 22.16 2.68 22.16 2.58 19.49 2.58  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.21 1.8 22.07 1.8 22.07 1.47 24.97 1.47 24.97 1.8 26.83 1.8 26.83 2.12 24.69 2.12 24.69 1.7 22.35 1.7 22.35 2.12 20.21 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.63 1.77 11.09 1.77 11.09 2.35 13.84 2.35 13.84 1.95 14.18 1.95 14.18 2.35 14.86 2.35 14.86 1.95 15.2 1.95 15.2 2.35 18.05 2.35 18.22 2.35 18.22 1.95 18.56 1.95 18.56 2.58 18.05 2.58 15.84 2.58 15.84 2.68 13.2 2.68 13.2 2.58 10.86 2.58 10.86 2.15 9.63 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.32 1.8 12.93 1.8 12.93 1.47 15.85 1.47 15.85 1.8 17.87 1.8 17.87 2.12 15.62 2.12 15.62 1.7 13.39 1.7 13.39 2.12 11.32 2.12  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.77 1.255 1.77 1.255 1.33 8.515 1.33 8.515 1.77 9.4 1.77 9.4 2.15 8.2 2.15 8.2 1.56 1.57 1.56 1.57 2.15 0.28 2.15  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.92 1.8 7.84 1.8 7.84 2.12 1.92 2.12  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.88075 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.12 2.82 21.91 2.82 21.91 2.92 25.05 2.92 25.05 2.82 27.965 2.82 27.965 2.53 28.195 2.53 28.195 3.38 27.965 3.38 27.965 3.05 25.3 3.05 25.3 3.24 21.66 3.24 21.66 3.05 19.12 3.05 19.12 3.38 18.81 3.38 18.81 3.05 18.05 3.05 16.34 3.05 16.34 3.24 12.7 3.24 12.7 3.05 6.66 3.05 6.66 3.24 4.955 3.24 4.955 3.38 4.725 3.38 4.725 3.24 3.02 3.24 3.02 3.05 0.525 3.05 0.525 3.38 0.295 3.38 0.295 2.53 0.525 2.53 0.525 2.82 4.725 2.82 4.725 2.53 4.955 2.53 4.955 2.82 12.95 2.82 12.95 2.92 16.09 2.92 16.09 2.82 18.05 2.82 18.81 2.82 18.81 0.99 27.01 0.99 27.01 1.22 19.12 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.28 2.77 3.28 2.77 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 12.11 3.62 12.11 3.285 12.45 3.285 12.45 3.62 16.59 3.62 16.59 3.285 16.93 3.285 16.93 3.62 18.05 3.62 21.07 3.62 21.07 3.285 21.41 3.285 21.41 3.62 25.55 3.62 25.55 3.285 25.89 3.285 25.89 3.62 28.36 3.62 28.56 3.62 28.56 4.22 28.36 4.22 18.05 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 28.56 -0.3 28.56 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.53 0.3 0.53 0.635 0.19 0.635 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.31 0.865 9.495 0.865 9.495 0.99 18.05 0.99 18.05 1.22 9.265 1.22 9.265 1.095 1.31 1.095  ;
        POLYGON 9.86 0.53 28.36 0.53 28.36 0.76 9.86 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_4
