# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.92 1.77 3.92 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.4295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 0.66 16.255 0.66 16.255 1.02 15.205 1.02 15.205 1.83 14.66 1.83  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.57 1.77 1.57 2.15 0.28 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.475 2.05 18.69 2.05 19.14 2.05 19.14 1.27 18.475 1.27 18.475 0.55 18.94 0.55 18.94 1.04 19.5 1.04 19.5 2.28 18.94 2.28 18.94 3.38 18.69 3.38 18.475 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.865 1.65 2.865 1.65 3.62 2.035 3.62 3.05 3.62 3.05 2.845 3.39 2.845 3.39 3.62 4.915 3.62 7.35 3.62 7.35 2.99 7.69 2.99 7.69 3.62 8.995 3.62 9.485 3.62 9.485 2.79 9.715 2.79 9.715 3.62 10.155 3.62 11.08 3.62 14.655 3.62 14.655 3.28 14.995 3.28 14.995 3.62 16.42 3.62 16.75 3.62 16.75 2.57 16.985 2.57 16.985 3.62 17.465 3.62 17.465 2.57 17.7 2.57 17.7 3.62 18.69 3.62 19.455 3.62 19.455 2.53 19.795 2.53 19.795 3.62 20.16 3.62 20.16 4.22 18.69 4.22 16.42 4.22 11.08 4.22 10.155 4.22 8.995 4.22 4.915 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.895 0.3 19.895 0.79 19.555 0.79 19.555 0.3 17.655 0.3 17.655 0.79 17.315 0.79 17.315 0.3 14.3 0.3 14.3 1.13 14.07 1.13 14.07 0.3 8.77 0.3 8.77 0.915 8.43 0.915 8.43 0.3 3.51 0.3 3.51 1.075 3.17 1.075 3.17 0.3 1.655 0.3 1.655 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.405 1.805 2.405 1.805 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.035 1.28 2.035 2.635 0.575 2.635 0.575 3.225 0.345 3.225  ;
        POLYGON 4.125 2.42 4.225 2.42 4.225 0.845 4.63 0.845 4.63 1.075 4.455 1.075 4.455 2.76 4.125 2.76  ;
        POLYGON 2.495 2.385 3.895 2.385 3.895 2.99 4.685 2.99 4.685 1.91 4.915 1.91 4.915 3.22 3.665 3.22 3.665 2.615 2.615 2.615 2.615 3.215 2.265 3.215 2.265 0.865 2.77 0.865 2.77 1.095 2.495 1.095  ;
        POLYGON 6.165 2.53 8.995 2.53 8.995 3.13 8.765 3.13 8.765 2.76 6.395 2.76 6.395 2.955 6.165 2.955  ;
        POLYGON 5.145 2.07 5.465 2.07 5.465 0.79 5.695 0.79 5.695 2.07 10.155 2.07 10.155 2.525 9.855 2.525 9.855 2.3 5.375 2.3 5.375 2.76 5.145 2.76  ;
        POLYGON 6.69 1.61 9.99 1.61 9.99 1 10.33 1 10.33 1.61 10.67 1.61 10.67 2.845 11.08 2.845 11.08 3.075 10.44 3.075 10.44 1.84 6.69 1.84  ;
        POLYGON 6.045 1.15 9 1.15 9 0.53 12.35 0.53 12.35 1.36 13.12 1.36 13.12 2.525 12.89 2.525 12.89 1.59 12.12 1.59 12.12 0.76 11.155 0.76 11.155 1.59 10.925 1.59 10.925 0.76 9.23 0.76 9.23 1.38 6.275 1.38 6.275 1.59 6.045 1.59  ;
        POLYGON 12.95 0.79 13.755 0.79 13.755 2.93 13.415 2.93 13.415 1.13 12.95 1.13  ;
        POLYGON 11.55 1 11.89 1 11.89 1.82 12.44 1.82 12.44 3.16 14.195 3.16 14.195 2.82 15.465 2.82 15.465 3.16 16.19 3.16 16.19 1.91 16.42 1.91 16.42 3.39 15.235 3.39 15.235 3.05 14.425 3.05 14.425 3.39 12.21 3.39 12.21 2.05 11.55 2.05  ;
        POLYGON 13.995 2.175 15.73 2.175 15.73 1.45 16.65 1.45 16.65 0.81 16.88 0.81 16.88 1.525 18.69 1.525 18.69 1.755 16.65 1.755 16.65 1.68 15.96 1.68 15.96 2.93 15.73 2.93 15.73 2.405 13.995 2.405  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
