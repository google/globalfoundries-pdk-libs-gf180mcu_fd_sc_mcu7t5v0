* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_2_3 net_2_3 A3 net_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_3 VSS A4 net_2_3 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_2 net_2_2 A4 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2_2 net_1 A3 net_2_2 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2_1 net_2_1 A3 net_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_1 VSS A4 net_2_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_0 net_2_0 A4 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_0 A3 net_2_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_3 net_0_3 A2 net_1_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_3 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_2 net_0_2 A1 ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_2 net_1 A2 net_0_2 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_1 net_0_1 A2 net_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_0 A1 ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_0 net_1 A2 net_0_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_6_3 ZN A3 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_7_3 VDD A4 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_7_2 ZN A4 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_6_2 VDD A3 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_6_1 ZN A3 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_7_1 VDD A4 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_7_0 ZN A4 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_6_0 VDD A3 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_5_3 ZN A2 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_4_3 VDD A1 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_4_2 ZN A1 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_5_2 VDD A2 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_5_1 ZN A2 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_4_1 VDD A1 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_4_0 ZN A1 VDD VNW pmos_5p0 W=8.45e-07 L=5e-07
M_i_5_0 VDD A2 ZN VNW pmos_5p0 W=8.45e-07 L=5e-07
.ENDS
