# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.685 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.105 1.535 10.785 1.535 10.785 1.21 11.235 1.21 12.755 1.21 12.755 1.59 11.235 1.59 11.065 1.59 11.065 1.765 10.105 1.765  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.865 1.77 2.71 1.77 2.71 3.27 2.33 3.27 2.33 2.15 1.865 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.29 1.77 1.59 1.77 1.59 2.15 0.29 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.924 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.7 2.33 17.57 2.33 18.01 2.33 18.01 1.535 14.82 1.535 14.82 0.705 15.05 0.705 15.05 1.265 17.06 1.265 17.06 0.705 17.29 0.705 17.29 1.265 18.39 1.265 18.39 2.71 17.57 2.71 16.99 2.71 16.99 3.195 16.76 3.195 16.76 2.71 14.975 2.71 14.975 3.195 14.7 3.195  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.28 3.62 6.28 2.605 6.51 2.605 6.51 3.62 9.69 3.62 9.69 2.92 9.92 2.92 9.92 3.62 11.635 3.62 11.635 2.76 11.865 2.76 11.865 3.62 13.7 3.62 13.7 3.04 13.93 3.04 13.93 3.62 15.74 3.62 15.74 3.04 15.97 3.04 15.97 3.62 17.57 3.62 17.78 3.62 17.78 3.045 18.01 3.045 18.01 3.62 19.04 3.62 19.04 4.22 17.57 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.41 0.3 18.41 0.805 18.18 0.805 18.18 0.3 16.17 0.3 16.17 0.805 15.94 0.805 15.94 0.3 13.93 0.3 13.93 0.805 13.7 0.805 13.7 0.3 10.05 0.3 10.05 0.845 9.82 0.845 9.82 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 0.995 1.31 0.995 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.765 0.53 0.765 0.53 1.225 1.885 1.225 1.885 0.765 2.77 0.765 2.77 0.995 2.115 0.995 2.115 1.46 0.19 1.46  ;
        POLYGON 3.46 1.445 3.69 1.445 3.69 1.87 4.935 1.87 4.935 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 5.205 2.33 5.205 1.34 7.08 1.34 7.08 1.575 5.435 1.575 5.435 2.56 4.04 2.56 4.04 3.125 3.81 3.125 3.81 2.56 3 2.56 3 0.765 3.89 0.765 3.89 0.995 3.23 0.995  ;
        POLYGON 7.915 0.53 9.075 0.53 9.075 0.76 8.275 0.76 8.275 1.805 8.93 1.805 8.93 2.85 8.645 2.85 8.645 2.035 7.915 2.035  ;
        POLYGON 9.175 1.075 10.28 1.075 10.28 0.53 11.235 0.53 11.235 0.76 10.51 0.76 10.51 1.305 9.415 1.305 9.415 1.995 10.945 1.995 10.945 2.85 10.715 2.85 10.715 2.225 9.175 2.225  ;
        POLYGON 5.685 1.805 7.32 1.805 7.32 0.78 7.55 0.78 7.55 3.16 9.165 3.16 9.165 2.455 10.43 2.455 10.43 3.16 11.175 3.16 11.175 1.995 13.075 1.995 13.075 1.965 13.415 1.965 13.415 2.225 11.405 2.225 11.405 3.39 10.2 3.39 10.2 2.69 9.395 2.69 9.395 3.39 7.32 3.39 7.32 2.035 5.685 2.035  ;
        POLYGON 12.68 2.455 13.7 2.455 13.7 1.535 13.105 1.535 13.105 0.76 11.595 0.76 11.595 0.53 13.335 0.53 13.335 1.265 13.93 1.265 13.93 1.825 17.57 1.825 17.57 2.095 13.93 2.095 13.93 2.685 12.91 2.685 12.91 3.265 12.68 3.265  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_4
