# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.65 1.8 8.415 1.8 8.415 2.12 1.65 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.795 1.325 8.04 1.325 8.04 1.22 9.42 1.22 9.42 2.255 9.06 2.255 9.06 1.56 0.795 1.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 0.865 1.365 0.865 1.365 0.53 1.595 0.53 1.595 0.865 3.605 0.865 3.605 0.53 3.835 0.53 3.835 0.865 5.845 0.865 5.845 0.53 6.075 0.53 6.075 0.865 7.5 0.865 7.5 0.53 8.41 0.53 8.41 0.76 7.73 0.76 7.73 1.095 0.43 1.095 0.43 2.35 7.195 2.35 7.195 3.38 6.965 3.38 6.965 2.7 5.65 2.7 5.65 2.585 3.87 2.585 3.87 2.7 2.715 2.7 2.715 3.38 2.485 3.38 2.485 2.7 1.17 2.7 1.17 2.585 0.13 2.585  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.24 3.62 0.24 2.815 0.58 2.815 0.58 3.62 4.67 3.62 4.67 2.815 5.01 2.815 5.01 3.62 9.1 3.62 9.1 2.815 9.44 2.815 9.44 3.62 10.08 3.62 10.08 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.5 0.3 9.5 0.635 9.14 0.635 9.14 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.54 0.3 0.54 0.635 0.18 0.635 0.18 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_4
