# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_64 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 35.84 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 6.245 3.62 6.245 2.49 6.475 2.49 6.475 3.62 8.485 3.62 8.485 2.49 8.715 2.49 8.715 3.62 10.725 3.62 10.725 2.49 10.955 2.49 10.955 3.62 12.965 3.62 12.965 2.49 13.195 2.49 13.195 3.62 15.205 3.62 15.205 2.49 15.435 2.49 15.435 3.62 17.445 3.62 17.445 2.49 17.675 2.49 17.675 3.62 19.685 3.62 19.685 2.49 19.915 2.49 19.915 3.62 21.925 3.62 21.925 2.49 22.155 2.49 22.155 3.62 24.165 3.62 24.165 2.49 24.395 2.49 24.395 3.62 26.405 3.62 26.405 2.49 26.635 2.49 26.635 3.62 28.645 3.62 28.645 2.49 28.875 2.49 28.875 3.62 30.885 3.62 30.885 2.49 31.115 2.49 31.115 3.62 33.125 3.62 33.125 2.49 33.355 2.49 33.355 3.62 35.365 3.62 35.365 2.49 35.595 2.49 35.595 3.62 35.84 3.62 35.84 4.22 35.595 4.22 33.355 4.22 31.115 4.22 28.875 4.22 26.635 4.22 24.395 4.22 22.155 4.22 19.915 4.22 17.675 4.22 15.435 4.22 13.195 4.22 10.955 4.22 8.715 4.22 6.475 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 35.84 -0.3 35.84 0.3 34.075 0.3 34.075 1.055 33.845 1.055 33.845 0.3 31.835 0.3 31.835 1.055 31.605 1.055 31.605 0.3 29.595 0.3 29.595 1.055 29.365 1.055 29.365 0.3 27.355 0.3 27.355 1.055 27.125 1.055 27.125 0.3 25.115 0.3 25.115 1.055 24.885 1.055 24.885 0.3 22.875 0.3 22.875 1.055 22.645 1.055 22.645 0.3 20.635 0.3 20.635 1.055 20.405 1.055 20.405 0.3 18.395 0.3 18.395 1.055 18.165 1.055 18.165 0.3 16.155 0.3 16.155 1.055 15.925 1.055 15.925 0.3 13.915 0.3 13.915 1.055 13.685 1.055 13.685 0.3 11.675 0.3 11.675 1.055 11.445 1.055 11.445 0.3 9.435 0.3 9.435 1.055 9.205 1.055 9.205 0.3 7.195 0.3 7.195 1.055 6.965 1.055 6.965 0.3 4.955 0.3 4.955 1.055 4.725 1.055 4.725 0.3 2.715 0.3 2.715 1.055 2.485 1.055 2.485 0.3 0.475 0.3 0.475 1.055 0.245 1.055 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
        POLYGON 4.725 1.325 6 1.325 6 1.555 4.955 1.555 4.955 3.39 4.725 3.39  ;
        POLYGON 5.21 1.96 6.245 1.96 6.245 0.53 6.475 0.53 6.475 2.19 5.21 2.19  ;
        POLYGON 6.965 1.325 8.24 1.325 8.24 1.555 7.195 1.555 7.195 3.39 6.965 3.39  ;
        POLYGON 7.45 1.96 8.485 1.96 8.485 0.53 8.715 0.53 8.715 2.19 7.45 2.19  ;
        POLYGON 9.205 1.325 10.48 1.325 10.48 1.555 9.435 1.555 9.435 3.39 9.205 3.39  ;
        POLYGON 9.69 1.96 10.725 1.96 10.725 0.53 10.955 0.53 10.955 2.19 9.69 2.19  ;
        POLYGON 11.445 1.325 12.72 1.325 12.72 1.555 11.675 1.555 11.675 3.39 11.445 3.39  ;
        POLYGON 11.93 1.96 12.965 1.96 12.965 0.53 13.195 0.53 13.195 2.19 11.93 2.19  ;
        POLYGON 13.685 1.325 14.96 1.325 14.96 1.555 13.915 1.555 13.915 3.39 13.685 3.39  ;
        POLYGON 14.17 1.96 15.205 1.96 15.205 0.53 15.435 0.53 15.435 2.19 14.17 2.19  ;
        POLYGON 15.925 1.325 17.2 1.325 17.2 1.555 16.155 1.555 16.155 3.39 15.925 3.39  ;
        POLYGON 16.41 1.96 17.445 1.96 17.445 0.53 17.675 0.53 17.675 2.19 16.41 2.19  ;
        POLYGON 18.165 1.325 19.44 1.325 19.44 1.555 18.395 1.555 18.395 3.39 18.165 3.39  ;
        POLYGON 18.65 1.96 19.685 1.96 19.685 0.53 19.915 0.53 19.915 2.19 18.65 2.19  ;
        POLYGON 20.405 1.325 21.68 1.325 21.68 1.555 20.635 1.555 20.635 3.39 20.405 3.39  ;
        POLYGON 20.89 1.96 21.925 1.96 21.925 0.53 22.155 0.53 22.155 2.19 20.89 2.19  ;
        POLYGON 22.645 1.325 23.92 1.325 23.92 1.555 22.875 1.555 22.875 3.39 22.645 3.39  ;
        POLYGON 23.13 1.96 24.165 1.96 24.165 0.53 24.395 0.53 24.395 2.19 23.13 2.19  ;
        POLYGON 24.885 1.325 26.16 1.325 26.16 1.555 25.115 1.555 25.115 3.39 24.885 3.39  ;
        POLYGON 25.37 1.96 26.405 1.96 26.405 0.53 26.635 0.53 26.635 2.19 25.37 2.19  ;
        POLYGON 27.125 1.325 28.4 1.325 28.4 1.555 27.355 1.555 27.355 3.39 27.125 3.39  ;
        POLYGON 27.61 1.96 28.645 1.96 28.645 0.53 28.875 0.53 28.875 2.19 27.61 2.19  ;
        POLYGON 29.365 1.325 30.64 1.325 30.64 1.555 29.595 1.555 29.595 3.39 29.365 3.39  ;
        POLYGON 29.85 1.96 30.885 1.96 30.885 0.53 31.115 0.53 31.115 2.19 29.85 2.19  ;
        POLYGON 31.605 1.325 32.88 1.325 32.88 1.555 31.835 1.555 31.835 3.39 31.605 3.39  ;
        POLYGON 32.09 1.96 33.125 1.96 33.125 0.53 33.355 0.53 33.355 2.19 32.09 2.19  ;
        POLYGON 33.845 1.325 35.12 1.325 35.12 1.555 34.075 1.555 34.075 3.39 33.845 3.39  ;
        POLYGON 34.33 1.96 35.365 1.96 35.365 0.53 35.595 0.53 35.595 2.19 34.33 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_64
