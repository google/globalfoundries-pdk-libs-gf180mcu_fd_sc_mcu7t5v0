# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 34.72 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.924 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.63 1.74 9.9 1.74 9.9 2.12 0.63 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.13 ;
    PORT
      LAYER METAL1 ;
        POLYGON 23.13 2.27 32.66 2.27 33.135 2.27 33.135 3.39 32.905 3.39 32.905 3 32.66 3 30.795 3 30.795 3.39 30.565 3.39 30.565 3 28.555 3 28.555 3.39 28.325 3.39 28.325 3 26.315 3 26.315 3.39 26.085 3.39 26.085 3 24.075 3 24.075 3.39 23.845 3.39 23.845 3 21.835 3 21.835 3.39 21.605 3.39 21.605 3 21.28 3 19.595 3 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 12.975 3 12.975 3.39 12.745 3.39 12.745 2.27 21.28 2.27 22.23 2.27 22.23 1.535 12.745 1.535 12.745 0.685 13.005 0.685 13.005 1.215 14.985 1.215 14.985 0.685 15.215 0.685 15.215 1.215 17.225 1.215 17.225 0.685 17.455 0.685 17.455 1.215 19.465 1.215 19.465 0.685 19.695 0.685 19.695 1.215 21.705 1.215 21.705 0.685 21.935 0.685 21.935 1.215 23.945 1.215 23.945 0.685 24.175 0.685 24.175 1.215 26.185 1.215 26.185 0.685 26.415 0.685 26.415 1.215 28.425 1.215 28.425 0.685 28.655 0.685 28.655 1.215 30.665 1.215 30.665 0.685 30.895 0.685 30.895 1.215 32.905 1.215 32.905 0.685 33.135 0.685 33.135 1.535 23.13 1.535  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.865 3.62 6.865 3.05 7.095 3.05 7.095 3.62 9.105 3.62 9.105 3.05 9.335 3.05 9.335 3.62 11.625 3.62 11.625 3.23 11.855 3.23 11.855 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.485 3.62 20.485 3.23 20.715 3.23 20.715 3.62 21.28 3.62 22.725 3.62 22.725 3.23 22.955 3.23 22.955 3.62 24.965 3.62 24.965 3.23 25.195 3.23 25.195 3.62 27.205 3.62 27.205 3.23 27.435 3.23 27.435 3.62 29.445 3.62 29.445 3.23 29.675 3.23 29.675 3.62 31.685 3.62 31.685 3.23 31.915 3.23 31.915 3.62 32.66 3.62 34.025 3.62 34.025 2.71 34.255 2.71 34.255 3.62 34.72 3.62 34.72 4.22 32.66 4.22 21.28 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 34.72 -0.3 34.72 0.3 34.255 0.3 34.255 1.05 34.025 1.05 34.025 0.3 32.07 0.3 32.07 0.985 31.73 0.985 31.73 0.3 29.83 0.3 29.83 0.985 29.49 0.985 29.49 0.3 27.59 0.3 27.59 0.985 27.25 0.985 27.25 0.3 25.35 0.3 25.35 0.985 25.01 0.985 25.01 0.3 23.11 0.3 23.11 0.985 22.77 0.985 22.77 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.675 0.3 11.675 1.04 11.445 1.04 11.445 0.3 9.435 0.3 9.435 1.04 9.205 1.04 9.205 0.3 7.195 0.3 7.195 1.04 6.965 1.04 6.965 0.3 4.955 0.3 4.955 1.04 4.725 1.04 4.725 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 2.53 10.325 2.53 10.325 1.505 1.365 1.505 1.365 0.685 1.595 0.685 1.595 1.27 3.605 1.27 3.605 0.685 3.835 0.685 3.835 1.27 5.845 1.27 5.845 0.685 6.075 0.685 6.075 1.27 8.085 1.27 8.085 0.685 8.315 0.685 8.315 1.27 10.325 1.27 10.325 0.685 10.555 0.685 10.555 1.765 21.28 1.765 21.28 1.995 10.555 1.995 10.555 3.39 10.325 3.39 10.325 2.82 8.215 2.82 8.215 3.39 7.985 3.39 7.985 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.595 2.76 1.595 3.39 1.365 3.39  ;
        POLYGON 23.86 1.765 32.66 1.765 32.66 1.995 23.86 1.995  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
