# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4685 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.89 1.77 4.03 1.77 4.03 2.15 2.89 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1415 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.09 1.77 15.285 1.77 15.285 2.15 14.09 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.765 1.59 1.765 1.59 2.13 0.28 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5972 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.05 2.06 21.605 2.06 22.01 2.06 22.01 1.315 20.045 1.315 20.045 0.55 20.28 0.55 20.28 1.085 22.01 1.085 22.01 0.55 22.535 0.55 22.535 3.38 21.67 3.38 21.67 2.29 21.605 2.29 20.28 2.29 20.28 3.38 20.05 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.09 3.62 3.24 3.62 3.24 2.845 3.58 2.845 3.58 3.62 5.115 3.62 7.675 3.62 7.675 3.445 8.015 3.445 8.015 3.62 10.275 3.62 10.275 3.005 10.615 3.005 10.615 3.62 12.315 3.62 14.295 3.62 14.295 3.005 14.635 3.005 14.635 3.62 15.6 3.62 16.705 3.62 16.705 2.53 16.935 2.53 16.935 3.62 18.75 3.62 18.75 2.53 18.98 2.53 18.98 3.62 21.17 3.62 21.17 2.53 21.4 2.53 21.4 3.62 21.605 3.62 23.41 3.62 23.41 2.53 23.64 2.53 23.64 3.62 24.08 3.62 24.08 4.22 21.605 4.22 15.6 4.22 12.315 4.22 5.115 4.22 2.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 23.64 0.3 23.64 0.89 23.41 0.89 23.41 0.3 21.455 0.3 21.455 0.835 21.115 0.835 21.115 0.3 19.08 0.3 19.08 0.89 18.85 0.89 18.85 0.3 16.895 0.3 16.895 0.835 16.555 0.835 16.555 0.3 7.795 0.3 7.795 1.075 7.455 1.075 7.455 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.36 1.86 2.36 1.86 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.09 1.28 2.09 2.595 0.575 2.595 0.575 3.225 0.345 3.225  ;
        POLYGON 4.27 0.79 4.61 0.79 4.61 2.93 4.27 2.93  ;
        POLYGON 2.62 2.38 4.04 2.38 4.04 3.16 4.885 3.16 4.885 1.93 5.115 1.93 5.115 3.39 3.81 3.39 3.81 2.615 2.615 2.615 2.615 3.225 2.385 3.225 2.385 0.81 2.715 0.81 2.715 1.15 2.62 1.15  ;
        POLYGON 5.345 0.79 5.675 0.79 5.675 1.765 8.235 1.765 8.235 1.995 5.575 1.995 5.575 2.985 5.345 2.985  ;
        POLYGON 6 1.305 8.11 1.305 8.11 0.53 11.04 0.53 11.04 1.615 10.81 1.615 10.81 0.76 8.34 0.76 8.34 1.535 6 1.535  ;
        POLYGON 7.015 2.225 9.035 2.225 9.035 2.08 9.875 2.08 9.875 0.99 10.215 0.99 10.215 2.08 11.645 2.08 11.645 2.78 11.305 2.78 11.305 2.31 9.375 2.31 9.375 2.93 9.035 2.93 9.035 2.455 7.015 2.455  ;
        POLYGON 6.115 2.24 6.455 2.24 6.455 2.985 8.5 2.985 8.5 3.16 9.685 3.16 9.685 2.54 11.075 2.54 11.075 3.065 12.315 3.065 12.315 3.295 10.845 3.295 10.845 2.775 9.915 2.775 9.915 3.39 8.27 3.39 8.27 3.215 6.115 3.215  ;
        POLYGON 13.86 2.54 15.6 2.54 15.6 2.885 15.37 2.885 15.37 2.775 13.86 2.775 13.86 2.845 13.63 2.845 13.63 1.22 12.555 1.22 12.555 0.99 14.495 0.99 14.495 1.22 13.86 1.22  ;
        POLYGON 11.27 0.79 11.93 0.79 11.93 0.53 16.11 0.53 16.11 1.395 17.335 1.395 17.335 1.63 15.88 1.63 15.88 0.76 12.16 0.76 12.16 2.55 12.895 2.55 12.895 2.78 11.93 2.78 11.93 1.13 11.27 1.13  ;
        POLYGON 15.755 1.86 17.73 1.86 17.73 0.55 17.96 0.55 17.96 1.555 21.605 1.555 21.605 1.785 17.96 1.785 17.96 3.38 17.73 3.38 17.73 2.105 15.755 2.105  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
