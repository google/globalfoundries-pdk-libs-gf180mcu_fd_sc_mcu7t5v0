# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.73 1.785 12.29 1.785 12.29 1.45 17.12 1.45 17.12 1.68 12.54 1.68 12.54 2.12 10.73 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.61 1.8 10.5 1.8 10.5 2.36 12.875 2.36 12.875 1.91 18.46 1.91 18.46 2.14 13.125 2.14 13.125 2.68 10.2 2.68 10.2 2.12 9.61 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.785 3.11 1.785 3.11 1.405 7.94 1.405 7.94 1.635 3.36 1.635 3.36 2.12 1.53 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.585 1.145 1.585 1.145 2.36 3.69 2.36 3.69 1.865 8.85 1.865 8.85 2.095 3.94 2.095 3.94 2.68 0.825 2.68  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.369 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 2.92 4.17 2.92 4.17 2.795 6.91 2.795 6.91 2.57 7.25 2.57 7.25 2.795 9.08 2.795 9.08 0.99 17.56 0.99 17.56 1.22 9.38 1.22 9.38 2.795 9.99 2.795 9.99 2.92 13.355 2.92 13.355 2.795 14.69 2.795 14.69 2.92 16.145 2.92 16.145 2.485 16.375 2.485 16.375 3.38 14.44 3.38 14.44 3.025 13.605 3.025 13.605 3.24 9.74 3.24 9.74 3.025 8.905 3.025 8.905 3.38 5.255 3.38 5.255 3.025 4.42 3.025 4.42 3.24 1.73 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.59 0.575 2.59 0.575 3.62 4.67 3.62 4.67 3.255 5.01 3.255 5.01 3.62 9.15 3.62 9.15 3.255 9.49 3.255 9.49 3.62 13.85 3.62 13.85 3.255 14.19 3.255 14.19 3.62 18.505 3.62 18.505 2.59 18.735 2.59 18.735 3.62 18.9 3.62 19.6 3.62 19.6 4.22 18.9 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.6 -0.3 19.6 0.3 8.37 0.3 8.37 0.715 8.03 0.715 8.03 0.3 6.13 0.3 6.13 0.715 5.79 0.715 5.79 0.3 3.89 0.3 3.89 0.715 3.55 0.715 3.55 0.3 1.65 0.3 1.65 0.715 1.31 0.715 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.55 0.53 0.55 0.53 0.945 2.43 0.945 2.43 0.55 2.77 0.55 2.77 0.945 4.67 0.945 4.67 0.55 5.01 0.55 5.01 0.945 6.91 0.945 6.91 0.55 7.25 0.55 7.25 0.945 8.61 0.945 8.61 0.53 18.9 0.53 18.9 0.76 8.84 0.76 8.84 1.175 0.19 1.175  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_4
