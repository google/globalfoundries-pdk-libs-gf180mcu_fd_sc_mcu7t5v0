# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.775 1.675 1.775 1.675 2.185 0.545 2.185  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.318 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.075 1.8 9.43 1.8 9.43 2.12 5.075 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.1496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.39 2.425 12.26 2.425 12.52 2.425 13.42 2.425 13.42 1.135 10.4 1.135 10.4 0.865 17.55 0.865 17.55 1.135 14.07 1.135 14.07 2.425 16.85 2.425 16.85 3.38 16.51 3.38 16.51 2.765 14.81 2.765 14.81 3.38 14.47 3.38 14.47 2.765 12.77 2.765 12.77 3.38 12.52 3.38 12.43 3.38 12.43 2.765 12.26 2.765 10.73 2.765 10.73 3.38 10.39 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.29 3.62 5.29 3.285 5.63 3.285 5.63 3.62 7.33 3.62 7.33 3.285 7.67 3.285 7.67 3.62 9.37 3.62 9.37 3.285 9.71 3.285 9.71 3.62 11.41 3.62 11.41 3.285 11.75 3.285 11.75 3.62 12.26 3.62 12.52 3.62 13.45 3.62 13.45 3.285 13.79 3.285 13.79 3.62 15.49 3.62 15.49 3.285 15.83 3.285 15.83 3.62 17.43 3.62 17.53 3.62 17.53 3.285 17.87 3.285 17.87 3.62 17.99 3.62 19.04 3.62 19.04 4.22 17.99 4.22 17.43 4.22 12.52 4.22 12.26 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.19 0.3 14.19 0.635 13.85 0.635 13.85 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.925 2.78 1.925 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.155 1.095 2.155 2.235 3.65 2.235 3.65 2.52 2.155 2.52 2.155 3.01 0.42 3.01  ;
        POLYGON 2.68 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.53 9.755 2.53 9.755 1.965 12.26 1.965 12.26 2.195 9.985 2.195 9.985 2.76 8.635 2.76 8.635 3.38 8.405 3.38 8.405 2.76 6.595 2.76 6.595 3.38 6.365 3.38 6.365 2.76 4.825 2.76 4.825 3.39 2.68 3.39  ;
        POLYGON 2.39 0.53 4.44 0.53 4.44 0.705 5.945 0.705 5.945 0.865 9.985 0.865 9.985 1.365 12.52 1.365 12.52 1.595 9.755 1.595 9.755 1.095 5.695 1.095 5.695 0.935 4.215 0.935 4.215 0.76 3.435 0.76 3.435 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 3.205 2.005 3.205 0.76 2.39 0.76  ;
        POLYGON 15.05 1.965 17.43 1.965 17.43 2.195 15.05 2.195  ;
        POLYGON 15.415 1.365 17.99 1.365 17.99 1.595 15.415 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_8
