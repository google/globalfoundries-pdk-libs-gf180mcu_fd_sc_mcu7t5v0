# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.01 1.24 2.325 1.24 2.325 0.55 2.7 0.55 2.7 1.59 2.01 1.59  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.78 1.82 2.95 1.82 2.95 1.27 3.21 1.27 3.21 1.82 4.045 1.82 4.045 2.795 3.49 2.795 3.49 2.12 0.78 2.12  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.39 1.8 7.39 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.86 2.11 14.37 2.11 14.67 2.11 14.67 1.39 11.825 1.39 11.825 0.545 12.055 0.545 12.055 1.16 14.065 1.16 14.065 0.545 14.295 0.545 14.295 1.16 15 1.16 15 2.34 14.46 2.34 14.46 3.38 14.37 3.38 13.965 3.38 13.965 2.34 12.22 2.34 12.22 3.38 11.86 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3 1.595 3 1.595 3.62 3.16 3.62 5.59 3.62 5.59 2.815 5.93 2.815 5.93 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 8.565 3.62 8.565 2.57 8.795 2.57 8.795 3.62 10.755 3.62 10.755 2.57 10.985 2.57 10.985 3.62 12.945 3.62 12.945 2.57 13.175 2.57 13.175 3.62 14.37 3.62 14.985 3.62 14.985 2.57 15.215 2.57 15.215 3.62 15.68 3.62 15.68 4.22 14.37 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 15.415 0.3 15.415 0.885 15.185 0.885 15.185 0.3 13.175 0.3 13.175 0.885 12.945 0.885 12.945 0.3 10.935 0.3 10.935 0.885 10.705 0.885 10.705 0.3 8.695 0.3 8.695 0.885 8.465 0.885 8.465 0.3 5.75 0.3 5.75 1.065 5.41 1.065 5.41 0.3 1.595 0.3 1.595 1.115 1.365 1.115 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.815 0.53 0.815 0.53 2.35 3.16 2.35 3.16 2.58 0.575 2.58 0.575 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 1.06 3.45 1.06 3.45 0.83 4.56 0.83 4.56 1.34 6.53 1.34 6.53 1.57 4.56 1.57 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.63 10.36 1.63 10.36 1.86 7.97 1.86 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 9.585 2.11 10.665 2.11 10.665 1.39 9.585 1.39 9.585 0.545 9.815 0.545 9.815 1.16 10.895 1.16 10.895 1.63 14.37 1.63 14.37 1.86 10.895 1.86 10.895 2.34 9.815 2.34 9.815 3.38 9.585 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_4
