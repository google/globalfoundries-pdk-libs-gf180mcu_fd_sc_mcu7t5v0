# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 1.765 6.155 1.765 6.155 2.15 0.64 2.15  ;
        POLYGON 7.8 1.765 13.31 1.765 13.31 2.15 7.8 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.0968 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.52 6.55 2.52 6.55 1.45 1.365 1.45 1.365 0.675 1.595 0.675 1.595 1.01 3.605 1.01 3.605 0.675 3.835 0.675 3.835 1.01 5.845 1.01 5.845 0.675 6.075 0.675 6.075 1.01 8.085 1.01 8.085 0.675 8.315 0.675 8.315 1.01 10.325 1.01 10.325 0.675 10.555 0.675 10.555 1.01 12.565 1.01 12.565 0.675 12.795 0.675 12.795 1.45 7.45 1.45 7.45 2.535 12.695 2.535 12.695 3.39 12.465 3.39 12.465 2.96 10.455 2.96 10.455 3.39 10.225 3.39 10.225 2.96 8.215 2.96 8.215 3.39 7.985 3.39 7.985 2.96 5.975 2.96 5.975 3.39 5.745 3.39 5.745 2.96 3.735 2.96 3.735 3.39 3.505 3.39 3.505 2.96 1.595 2.96 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.68 0.475 2.68 0.475 3.62 2.385 3.62 2.385 3.21 2.615 3.21 2.615 3.62 4.625 3.62 4.625 3.21 4.855 3.21 4.855 3.62 6.865 3.62 6.865 3.21 7.095 3.21 7.095 3.62 9.105 3.62 9.105 3.21 9.335 3.21 9.335 3.62 11.345 3.62 11.345 3.21 11.575 3.21 11.575 3.62 13.585 3.62 13.585 2.68 13.815 2.68 13.815 3.62 14.56 3.62 14.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.915 0.3 13.915 1.015 13.685 1.015 13.685 0.3 11.675 0.3 11.675 0.69 11.445 0.69 11.445 0.3 9.435 0.3 9.435 0.69 9.205 0.69 9.205 0.3 7.195 0.3 7.195 0.69 6.965 0.69 6.965 0.3 4.955 0.3 4.955 0.69 4.725 0.69 4.725 0.3 2.715 0.3 2.715 0.69 2.485 0.69 2.485 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_12
