# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.88 1.265 4.36 1.265 4.36 1.535 1.88 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 1.6 1.105 1.6 1.105 2.225 3.41 2.225 3.645 2.225 3.645 1.82 4.615 1.82 4.615 1.56 5.36 1.56 5.36 1.79 4.895 1.79 4.895 2.095 3.875 2.095 3.875 2.455 3.41 2.455 2.1 2.455 2.1 2.71 0.865 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.4355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.91 1.82 9.555 1.82 10.6 1.82 10.6 2.115 9.555 2.115 7.91 2.115  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.025 2.36 17.225 2.36 17.48 2.36 17.48 1.56 13.025 1.56 13.025 0.6 13.335 0.6 13.335 1.24 15.265 1.24 15.265 0.6 15.575 0.6 15.575 1.24 17.505 1.24 17.505 0.6 17.815 0.6 17.815 3.325 17.37 3.325 17.37 2.68 17.225 2.68 15.69 2.68 15.69 3.315 15.265 3.315 15.265 2.68 13.505 2.68 13.505 3.315 13.025 3.315  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.33 3.62 2.33 2.685 2.67 2.685 2.67 3.62 3.41 3.62 5.875 3.62 6.365 3.62 6.365 2.485 6.595 2.485 6.595 3.62 8.57 3.62 8.57 2.805 8.91 2.805 8.91 3.62 12.23 3.62 12.23 3.285 12.57 3.285 12.57 3.62 14.225 3.62 14.225 2.94 14.455 2.94 14.455 3.62 16.415 3.62 16.415 2.94 16.645 2.94 16.645 3.62 17.225 3.62 18.48 3.62 18.48 4.22 17.225 4.22 5.875 4.22 3.41 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.695 0.3 16.695 0.84 16.465 0.84 16.465 0.3 14.455 0.3 14.455 0.85 14.225 0.85 14.225 0.3 8.69 0.3 8.69 0.775 8.35 0.775 8.35 0.3 5.93 0.3 5.93 0.76 5.59 0.76 5.59 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.085 1.12 1.58 1.12 1.58 1.765 3.41 1.765 3.41 1.995 1.35 1.995 1.35 1.355 0.575 1.355 0.575 2.98 0.345 2.98 0.345 1.12 0.835 1.12 0.835 0.53 1.65 0.53 1.65 0.76 1.085 0.76  ;
        POLYGON 3.55 2.685 3.89 2.685 3.89 3.16 5.645 3.16 5.645 2.61 5.875 2.61 5.875 3.39 3.55 3.39  ;
        POLYGON 6.31 0.53 7.615 0.53 7.615 1.35 9.555 1.35 9.555 1.585 7.615 1.585 7.615 2.845 7.385 2.845 7.385 0.765 6.31 0.765  ;
        POLYGON 4.57 2.685 5.14 2.685 5.14 2.025 5.705 2.025 5.705 1.305 5.035 1.305 5.035 0.76 3.55 0.76 3.55 0.53 5.265 0.53 5.265 1.075 7.115 1.075 7.115 3.14 7.97 3.14 7.97 2.345 11.765 2.345 11.765 1.695 11.995 1.695 11.995 2.575 8.205 2.575 8.205 3.39 6.885 3.39 6.885 1.305 5.935 1.305 5.935 2.26 5.37 2.26 5.37 2.915 4.57 2.915  ;
        POLYGON 9.56 0.53 12.68 0.53 12.68 0.76 9.56 0.76  ;
        POLYGON 9.635 2.815 12.345 2.815 12.345 1.22 10.98 1.22 10.98 0.99 12.575 0.99 12.575 1.825 17.225 1.825 17.225 2.095 12.575 2.095 12.575 3.05 9.635 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_4
