# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4635 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7115 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5259 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.49 2.245 17.91 2.245 18.57 2.245 18.57 1.555 16.49 1.555 16.49 0.99 16.83 0.99 16.83 1.325 19.17 1.325 19.17 0.99 19.51 0.99 19.51 2.93 18.87 2.93 18.87 2.595 17.91 2.595 16.84 2.595 16.84 2.93 16.49 2.93  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.44 3.62 1.44 2.93 1.78 2.93 1.78 3.62 2.165 3.62 3.18 3.62 3.18 3.005 3.52 3.005 3.52 3.62 6.355 3.62 7.705 3.62 7.705 2.7 8.045 2.7 8.045 3.62 9.38 3.62 12.85 3.62 12.85 3.28 13.19 3.28 13.19 3.62 15.25 3.62 15.25 2.815 15.59 2.815 15.59 3.62 17.73 3.62 17.73 3.285 18.07 3.285 18.07 3.62 20.13 3.62 20.51 3.62 20.51 2.815 20.85 2.815 20.85 3.62 21.28 3.62 21.28 4.22 20.13 4.22 9.38 4.22 6.355 4.22 2.165 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.795 0.3 20.795 0.765 20.565 0.765 20.565 0.3 18.17 0.3 18.17 0.635 17.83 0.635 17.83 0.3 15.435 0.3 15.435 0.69 15.205 0.69 15.205 0.3 13.19 0.3 13.19 0.635 12.85 0.635 12.85 0.3 8.04 0.3 8.04 0.81 7.7 0.81 7.7 0.3 3.62 0.3 3.62 1.075 3.28 1.075 3.28 0.3 1.78 0.3 1.78 0.915 1.44 0.915 1.44 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.475 2.36 1.935 2.36 1.935 1.375 0.375 1.375 0.375 0.735 0.605 0.735 0.605 1.145 2.165 1.145 2.165 2.59 0.705 2.59 0.705 3.225 0.475 3.225  ;
        POLYGON 4.42 2.645 5.055 2.645 5.055 1.075 4.4 1.075 4.4 0.845 5.29 0.845 5.29 2.875 4.42 2.875  ;
        POLYGON 2.515 0.735 2.845 0.735 2.845 2.48 4.06 2.48 4.06 3.16 6.355 3.16 6.355 3.39 3.83 3.39 3.83 2.71 2.845 2.71 2.845 3.225 2.515 3.225  ;
        POLYGON 5.575 0.79 5.805 0.79 5.805 1.82 6.55 1.82 6.55 1.5 8.7 1.5 8.7 1.73 6.78 1.73 6.78 2.05 5.915 2.05 5.915 2.795 5.575 2.795  ;
        POLYGON 7.095 2.05 9.04 2.05 9.04 0.99 9.38 0.99 9.38 2.93 9.04 2.93 9.04 2.39 7.095 2.39  ;
        POLYGON 6.09 1.04 8.33 1.04 8.33 0.53 11.51 0.53 11.51 2.04 11.17 2.04 11.17 0.76 8.56 0.76 8.56 1.27 6.32 1.27 6.32 1.59 6.09 1.59  ;
        POLYGON 10.16 0.99 10.5 0.99 10.5 2.355 13.43 2.355 13.43 2.105 13.77 2.105 13.77 2.585 10.5 2.585 10.5 2.93 10.16 2.93  ;
        POLYGON 12.41 1.495 14.15 1.495 14.15 0.99 14.49 0.99 14.49 1.785 17.91 1.785 17.91 2.015 14.43 2.015 14.43 2.795 14.09 2.795 14.09 1.73 12.41 1.73  ;
        POLYGON 11.79 2.815 13.73 2.815 13.73 3.025 14.79 3.025 14.79 2.295 16.055 2.295 16.055 3.16 17.27 3.16 17.27 2.825 18.53 2.825 18.53 3.16 19.9 3.16 19.9 0.76 18.63 0.76 18.63 1.095 17.37 1.095 17.37 0.76 15.895 0.76 15.895 1.15 14.745 1.15 14.745 0.76 13.65 0.76 13.65 1.095 11.745 1.095 11.745 0.675 11.975 0.675 11.975 0.865 13.42 0.865 13.42 0.53 14.975 0.53 14.975 0.92 15.665 0.92 15.665 0.53 17.6 0.53 17.6 0.865 18.4 0.865 18.4 0.53 20.13 0.53 20.13 3.39 18.3 3.39 18.3 3.055 17.5 3.055 17.5 3.39 15.825 3.39 15.825 2.525 15.02 2.525 15.02 3.255 13.5 3.255 13.5 3.05 11.79 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_4
