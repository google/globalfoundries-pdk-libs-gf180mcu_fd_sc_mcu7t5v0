# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.24 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.05 1.265 4.535 1.265 4.535 1.535 2.05 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.075 1.49 1.305 1.49 1.305 2.225 3.56 2.225 3.835 2.225 3.835 1.765 4.8 1.765 4.8 1.485 5.695 1.485 5.695 1.72 5.095 1.72 5.095 2.095 4.065 2.095 4.065 2.455 3.56 2.455 2.275 2.455 2.275 2.66 1.075 2.66  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.115 1.825 9.61 1.825 10.71 1.825 10.71 2.095 9.61 2.095 8.115 2.095  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7952 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.29 2.36 15.21 2.36 15.46 2.36 15.46 1.56 13.29 1.56 13.29 0.655 13.52 0.655 13.52 1.24 15.53 1.24 15.53 0.655 15.76 0.655 15.76 3.36 15.24 3.36 15.24 2.68 15.21 2.68 13.52 2.68 13.52 3.36 13.29 3.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.725 3.62 2.725 2.735 3.065 2.735 3.065 3.62 3.56 3.62 6.07 3.62 6.525 3.62 6.525 2.68 6.81 2.68 6.81 3.62 8.775 3.62 8.775 2.795 9.135 2.795 9.135 3.62 11.99 3.62 11.99 3.28 12.355 3.28 12.355 3.62 14.31 3.62 14.31 3.015 14.54 3.015 14.54 3.62 15.21 3.62 16.24 3.62 16.24 4.22 15.21 4.22 6.07 4.22 3.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 16.24 -0.3 16.24 0.3 14.64 0.3 14.64 0.905 14.41 0.905 14.41 0.3 8.88 0.3 8.88 0.76 8.535 0.76 8.535 0.3 6.095 0.3 6.095 0.76 5.755 0.76 5.755 0.3 2.935 0.3 2.935 0.775 2.595 0.775 2.595 0.3 0.695 0.3 0.695 0.76 0.355 0.76 0.355 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.51 0.99 1.475 0.99 1.475 0.53 1.815 0.53 1.815 1.765 3.56 1.765 3.56 1.995 1.535 1.995 1.535 1.22 0.74 1.22 0.74 3.03 0.51 3.03  ;
        POLYGON 3.735 2.735 4.095 2.735 4.095 3.16 5.785 3.16 5.785 2.68 6.07 2.68 6.07 3.39 3.735 3.39  ;
        POLYGON 6.485 0.53 7.885 0.53 7.885 0.99 9.61 0.99 9.61 1.555 9.27 1.555 9.27 1.22 7.885 1.22 7.885 2.78 7.545 2.78 7.545 0.76 6.485 0.76  ;
        POLYGON 4.72 2.605 5.325 2.605 5.325 1.99 7.01 1.99 7.01 1.22 5.24 1.22 5.24 0.76 3.625 0.76 3.625 0.53 5.47 0.53 5.47 0.99 7.27 0.99 7.27 3.01 8.16 3.01 8.16 2.33 11.105 2.33 11.105 1.67 11.76 1.67 11.76 1.9 11.335 1.9 11.335 2.565 8.445 2.565 8.445 3.24 7.04 3.24 7.04 2.22 5.555 2.22 5.555 2.835 4.72 2.835  ;
        POLYGON 9.795 0.53 12.865 0.53 12.865 0.76 9.795 0.76  ;
        POLYGON 9.75 2.815 12.125 2.815 12.125 1.22 11.17 1.22 11.17 0.99 12.355 0.99 12.355 1.825 15.21 1.825 15.21 2.095 12.355 2.095 12.355 3.05 9.75 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_2
