# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 32.48 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.5485 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.69 1.77 12.79 1.77 12.79 2.15 5.69 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.2992 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.95 2.505 21.92 2.505 22.23 2.505 22.23 1.095 14.97 1.095 14.97 0.865 30.99 0.865 30.99 1.095 23.13 1.095 23.13 2.505 29.57 2.505 29.57 3.38 29.23 3.38 29.23 3.055 27.53 3.055 27.53 3.38 27.19 3.38 27.19 3.055 25.49 3.055 25.49 3.38 25.15 3.38 25.15 3.055 23.45 3.055 23.45 3.38 23.13 3.38 23.13 3.055 21.92 3.055 21.41 3.055 21.41 3.38 21.07 3.38 21.07 3.055 19.37 3.055 19.37 3.38 19.03 3.38 19.03 3.055 17.33 3.055 17.33 3.38 16.99 3.38 16.99 3.055 15.29 3.055 15.29 3.38 14.95 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.29 3.62 5.29 3.04 5.63 3.04 5.63 3.62 7.33 3.62 7.33 3.04 7.67 3.04 7.67 3.62 9.37 3.62 9.37 3.04 9.71 3.04 9.71 3.62 11.71 3.62 11.71 3.04 12.05 3.04 12.05 3.62 13.93 3.62 13.93 2.53 14.27 2.53 14.27 3.62 15.97 3.62 15.97 3.285 16.31 3.285 16.31 3.62 18.01 3.62 18.01 3.285 18.35 3.285 18.35 3.62 20.05 3.62 20.05 3.285 20.39 3.285 20.39 3.62 21.92 3.62 22.09 3.62 22.09 3.285 22.43 3.285 22.43 3.62 24.13 3.62 24.13 3.285 24.47 3.285 24.47 3.62 26.17 3.62 26.17 3.285 26.51 3.285 26.51 3.62 28.21 3.62 28.21 3.285 28.55 3.285 28.55 3.62 30.08 3.62 30.305 3.62 30.305 2.53 30.535 2.53 30.535 3.62 31.52 3.62 32.48 3.62 32.48 4.22 31.52 4.22 30.08 4.22 21.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 32.48 -0.3 32.48 0.3 32.055 0.3 32.055 0.9 31.825 0.9 31.825 0.3 29.87 0.3 29.87 0.635 29.53 0.635 29.53 0.3 27.63 0.3 27.63 0.635 27.29 0.635 27.29 0.3 25.39 0.3 25.39 0.635 25.05 0.635 25.05 0.3 23.15 0.3 23.15 0.635 22.81 0.635 22.81 0.3 20.91 0.3 20.91 0.635 20.57 0.635 20.57 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.21 0.3 14.21 0.635 13.835 0.635 13.835 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.42 2.78 1.895 2.78 1.895 1.325 0.19 1.325 0.19 0.865 0.53 0.865 0.53 1.095 2.125 1.095 2.125 2.235 3.65 2.235 3.65 2.52 2.125 2.52 2.125 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 6.35 0.705 6.35 0.865 13.64 0.865 13.64 1.36 21.45 1.36 21.45 1.59 13.35 1.59 13.35 1.095 6.01 1.095 6.01 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.73 3.16 4.83 3.16 4.83 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 5.06 1.315 5.06 2.53 13.27 2.53 13.27 2 21.92 2 21.92 2.23 13.615 2.23 13.615 2.76 13.13 2.76 13.13 3.38 12.79 3.38 12.79 2.76 10.885 2.76 10.885 3.38 10.545 3.38 10.545 2.76 8.69 2.76 8.69 3.38 8.35 3.38 8.35 2.76 6.65 2.76 6.65 3.38 6.31 3.38 6.31 2.76 5.06 2.76 5.06 3.39 2.73 3.39  ;
        POLYGON 23.63 2 30.08 2 30.08 2.23 23.63 2.23  ;
        POLYGON 23.49 1.36 31.52 1.36 31.52 1.59 23.49 1.59  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_16
