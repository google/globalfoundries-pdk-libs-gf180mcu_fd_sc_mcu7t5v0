# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.16 1.77 8.82 1.77 8.82 2.365 11.34 2.365 11.34 1.77 12.59 1.77 12.59 2.15 11.57 2.15 11.57 2.595 8.55 2.595 8.55 2.15 8.16 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.05 1.8 11.11 1.8 11.11 2.12 9.05 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.53 1.8 4.71 1.8 4.71 2.12 1.53 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.625 1.16 1.69 1.16 1.69 1.34 4.455 1.34 4.455 1.57 1 1.57 1 2.275 0.625 2.275  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.105 1.8 6.865 1.8 7.33 1.8 7.33 2.12 6.865 2.12 5.105 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.382 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.915 2.825 12.58 2.825 12.58 3.26 10.525 3.26 10.525 3.055 9.54 3.055 9.54 3.26 7.56 3.26 7.56 2.68 6.865 2.68 5.775 2.68 5.775 3.11 5.545 3.11 5.545 2.68 2.715 2.68 2.715 3.375 2.485 3.375 2.485 2.36 6.865 2.36 7.56 2.36 7.56 0.99 11.33 0.99 11.33 1.22 7.915 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.69 0.475 2.69 0.475 3.62 4.67 3.62 4.67 3.09 5.01 3.09 5.01 3.62 6.51 3.62 6.51 3.09 6.85 3.09 6.85 3.62 6.865 3.62 9.87 3.62 9.87 3.285 10.21 3.285 10.21 3.62 12.68 3.62 12.88 3.62 12.88 4.22 12.68 4.22 6.865 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 5.01 0.3 5.01 0.635 4.665 0.635 4.665 0.3 2.77 0.3 2.77 0.635 2.425 0.635 2.425 0.3 0.53 0.3 0.53 0.635 0.185 0.635 0.185 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.26 0.55 2.17 0.55 2.17 0.865 5.11 0.865 5.11 0.99 6.865 0.99 6.865 1.22 4.86 1.22 4.86 1.095 1.94 1.095 1.94 0.78 1.26 0.78  ;
        POLYGON 5.38 0.53 12.68 0.53 12.68 0.76 5.38 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_2
