* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24 net_7 net_9 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55 net_6 net_8 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27 net_17 net_14 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63 net_16 net_15 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22 net_13 net_11 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93 net_12 net_10 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_20 net_30 net_26 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_59 net_25 net_20 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_135 net_23 net_28 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_90 net_33 net_18 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27_139 net_31 net_29 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63_82 net_32 net_24 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22_30 net_22 net_27 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93_110 net_19 net_21 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33 VDD net_7 net_9 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23 VDD net_6 net_8 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94 VDD net_17 net_14 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87 VDD net_16 net_15 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95 VDD net_13 net_11 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23 VDD net_12 net_10 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_95 VDD net_30 net_26 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_188 VDD net_25 net_20 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_98 VDD net_23 net_28 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_16 VDD net_33 net_18 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94_91 VDD net_31 net_29 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87_65 VDD net_32 net_24 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95_109 VDD net_22 net_27 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23_99 VDD net_19 net_21 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS
