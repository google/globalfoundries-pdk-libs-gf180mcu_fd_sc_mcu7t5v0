# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.18 1.8 14.73 1.8 14.73 2.12 11.18 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.445 1.71 10.16 1.71 10.16 1.24 13.78 1.24 13.78 0.53 17.05 0.53 17.05 2.235 16.82 2.235 16.82 0.76 14.01 0.76 14.01 1.56 10.52 1.56 10.52 2.14 9.445 2.14  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.64 1.8 7.24 1.8 7.24 2.13 1.64 2.13  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.23 3.375 1.23 3.375 1.325 8.12 1.325 8.12 1.56 1.02 1.56 1.02 2.225 0.62 2.225  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.215 2.67 15.05 2.67 15.05 0.99 15.58 0.99 15.58 2.67 16.67 2.67 16.67 2.91 8.985 2.91 8.985 1.095 3.765 1.095 3.765 0.8 2.225 0.8 2.225 0.57 3.995 0.57 3.995 0.865 6.365 0.865 6.365 0.57 6.595 0.57 6.595 0.865 8.985 0.865 8.985 0.53 11.18 0.53 11.18 1 9.215 1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 3.01 1.55 3.01 1.55 3.62 3.25 3.62 3.25 3.01 3.59 3.01 3.59 3.62 5.29 3.62 5.29 3.01 5.63 3.01 5.63 3.62 7.33 3.62 7.33 3.01 7.67 3.01 7.67 3.62 17.65 3.62 17.92 3.62 17.92 4.22 17.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 17.595 0.3 17.595 0.73 17.365 0.73 17.365 0.3 13.075 0.3 13.075 0.73 12.845 0.73 12.845 0.3 8.69 0.3 8.69 0.635 8.35 0.635 8.35 0.3 4.61 0.3 4.61 0.635 4.27 0.635 4.27 0.3 0.475 0.3 0.475 0.695 0.245 0.695 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 2.485 8.69 2.485 8.69 3.16 17.31 3.16 17.31 2.485 17.65 2.485 17.65 3.39 8.35 3.39 8.35 2.715 6.65 2.715 6.65 3.39 6.31 3.39 6.31 2.715 4.61 2.715 4.61 3.39 4.27 3.39 4.27 2.715 2.57 2.715 2.57 3.39 2.23 3.39 2.23 2.715 0.53 2.715 0.53 3.39 0.19 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_4
