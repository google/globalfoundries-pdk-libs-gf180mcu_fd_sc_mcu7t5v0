# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.84 1.73 1.56 1.73 1.56 3.38 1.22 3.38 1.22 2.14 0.84 2.14  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 1.61 2.14 1.61 2.14 3.38 1.79 3.38  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.9 1.61 3.26 1.61 3.26 3.38 2.9 3.38  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.84 2.38 5.515 2.38 5.745 2.38 5.745 1.535 4.87 1.535 4.87 0.53 5.49 0.53 5.49 1.265 6.04 1.265 6.04 2.655 5.515 2.655 5.46 2.655 5.46 3.38 4.84 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 3.715 3.62 3.715 2.53 3.945 2.53 3.945 3.62 5.515 3.62 5.925 3.62 5.925 2.935 6.155 2.935 6.155 3.62 6.72 3.62 6.72 4.22 5.515 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 6.255 0.3 6.255 0.92 6.025 0.92 6.025 0.3 3.835 0.3 3.835 0.895 3.605 0.895 3.605 0.3 1.595 0.3 1.595 0.895 1.365 0.895 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.53 0.475 0.53 0.475 1.125 2.485 1.125 2.485 0.53 2.715 0.53 2.715 1.125 4.19 1.125 4.19 1.765 5.515 1.765 5.515 1.995 3.96 1.995 3.96 1.36 0.575 1.36 0.575 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_2
