# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.19 1.035 1.19 1.035 1.735 1.97 1.735 1.97 2.12 1.035 2.12 1.035 2.875 0.705 2.875  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.006 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 2.33 2.36 2.33 1.505 1.365 1.505 1.365 0.68 1.595 0.68 1.595 1.27 2.71 1.27 2.71 2.735 1.495 2.735 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 3.36 3.62 3.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_2
