# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.76 1.62 1.76 1.62 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.475 1.79 6.07 1.79 6.07 2.135 4.475 2.135  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.08 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 2.425 9.95 2.425 10.125 2.425 10.73 2.425 10.73 1.1 9.4 1.1 9.4 0.715 9.63 0.715 9.63 0.865 11.64 0.865 11.64 0.71 11.87 0.71 11.87 1.1 11.11 1.1 11.11 2.425 11.42 2.425 11.42 3.38 11.19 3.38 11.19 2.66 10.125 2.66 9.95 2.66 9.41 2.66 9.41 3.38 9.11 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.455 3.62 1.455 3.285 1.795 3.285 1.795 3.62 5.985 3.62 5.985 3.285 6.325 3.285 6.325 3.62 8.075 3.62 8.075 2.815 8.415 2.815 8.415 3.62 9.95 3.62 10.125 3.62 10.17 3.62 10.17 3.02 10.4 3.02 10.4 3.62 12.21 3.62 12.21 2.565 12.44 2.565 12.44 3.62 13.44 3.62 13.44 4.22 10.125 4.22 9.95 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 12.99 0.3 12.99 1.06 12.76 1.06 12.76 0.3 10.805 0.3 10.805 0.635 10.465 0.635 10.465 0.3 8.565 0.3 8.565 0.635 8.225 0.635 8.225 0.3 6.325 0.3 6.325 0.635 5.985 0.635 5.985 0.3 1.595 0.3 1.595 0.76 1.365 0.76 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.49 2.51 1.87 2.51 1.87 1.225 0.245 1.225 0.245 0.67 0.475 0.67 0.475 0.99 2.1 0.99 2.1 2.085 3.26 2.085 3.26 2.32 2.1 2.32 2.1 2.74 0.72 2.74 0.72 3.38 0.49 3.38  ;
        POLYGON 4.89 2.365 6.6 2.365 6.6 1.56 4.935 1.56 4.935 1.22 4.515 1.22 4.515 0.99 5.165 0.99 5.165 1.325 6.83 1.325 6.83 1.73 7.94 1.73 7.94 2.125 6.83 2.125 6.83 2.595 5.12 2.595 5.12 2.89 4.89 2.89  ;
        POLYGON 2.475 3.125 4.01 3.125 4.01 1.345 3.76 1.345 3.76 0.99 4.24 0.99 4.24 3.12 5.395 3.12 5.395 2.825 7.11 2.825 7.11 2.355 8.335 2.355 8.335 1.96 9.95 1.96 9.95 2.195 8.565 2.195 8.565 2.585 7.34 2.585 7.34 3.38 7.11 3.38 7.11 3.055 5.625 3.055 5.625 3.355 2.475 3.355  ;
        POLYGON 2.485 0.53 5.625 0.53 5.625 0.865 8.565 0.865 8.565 1.365 10.125 1.365 10.125 1.595 8.335 1.595 8.335 1.095 5.395 1.095 5.395 0.76 3.205 0.76 3.205 1.575 3.78 1.575 3.78 2.89 3.545 2.89 3.545 1.805 2.975 1.805 2.975 0.885 2.485 0.885  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_4
