# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 1.75 1.79 1.75 1.79 1.16 2.13 1.16 2.13 2.15 1.23 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 1.47 3.81 1.47 3.81 3.32 3.47 3.32  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 1.47 4.935 1.47 4.935 3.32 4.59 3.32  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.054 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.16 1 1.16 1 3.32 0.705 3.32  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.33 2.38 2.36 2.38 2.36 0.99 4.33 0.99 5.165 0.99 5.165 0.605 5.395 0.605 5.395 1.22 4.33 1.22 2.68 1.22 2.68 2.68 1.67 2.68 1.67 3.38 1.33 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 4.33 3.62 5.165 3.62 5.165 2.53 5.395 2.53 5.395 3.62 6.16 3.62 6.16 4.22 4.33 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 0.475 0.3 0.475 0.945 0.245 0.945 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 0.53 4.33 0.53 4.33 0.76 1.31 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_1
