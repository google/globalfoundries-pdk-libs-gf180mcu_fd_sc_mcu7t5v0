# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 8.96 3.62 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_16
