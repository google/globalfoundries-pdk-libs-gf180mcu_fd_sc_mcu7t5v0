# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.04 1.525 4.36 1.525 4.36 3.32 4.04 3.32  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.16 1.77 6.04 1.77 6.04 2.14 5.48 2.14 5.48 3.32 5.16 3.32  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.28 1.77 6.57 1.77 7.87 1.77 7.87 2.14 6.6 2.14 6.6 3.32 6.57 3.32 6.28 3.32  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.92 1.525 3.24 1.525 3.24 3.32 2.92 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.8 1.525 2.12 1.525 2.12 3.32 1.8 3.32  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 1.525 1 1.525 1 3.32 0.705 3.32  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.8719 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.49 0.99 6.57 0.99 7.405 0.99 7.405 0.555 7.635 0.555 7.635 1.22 6.57 1.22 3.79 1.22 3.79 3.38 3.49 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 6.57 3.62 7.305 3.62 7.305 2.53 7.535 2.53 7.535 3.62 8.4 3.62 8.4 4.22 6.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 2.715 0.3 2.715 0.815 2.485 0.815 2.485 0.3 0.475 0.3 0.475 0.815 0.245 0.815 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 0.53 1.595 0.53 1.595 1.045 2.945 1.045 2.945 0.53 6.57 0.53 6.57 0.76 3.175 0.76 3.175 1.275 1.365 1.275  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_1
