# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.8 1.45 13.38 1.45 13.38 1.16 14.42 1.16 14.44 1.16 14.44 2.38 14.42 2.38 14.12 2.38 14.12 1.68 9.8 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.48 1.78 9.52 1.78 9.52 1.91 12.54 1.91 12.54 2.14 8.48 2.14  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.44 1.78 8.23 1.78 8.23 2.37 13.435 2.37 13.435 1.91 13.775 1.91 13.775 2.68 8 2.68 8 2.14 7.44 2.14  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.89 1.8 4.95 1.8 4.95 2.12 2.89 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.51 1.77 2.41 1.77 2.41 1.325 5.48 1.325 5.48 2.15 5.18 2.15 5.18 1.555 2.66 1.555 2.66 2.15 1.51 2.15  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.8 1.145 1.8 1.145 2.38 5.72 2.38 5.72 1.8 6.6 1.8 6.6 2.12 6.06 2.12 6.06 2.68 0.825 2.68 0.825 2.12 0.28 2.12  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.8038 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.75 2.92 6.41 2.92 6.41 2.825 6.85 2.825 6.85 0.99 13.07 0.99 13.07 1.22 7.15 1.22 7.15 2.825 7.75 2.825 7.75 2.92 11.215 2.92 11.215 3.24 7.5 3.24 7.5 3.055 6.66 3.055 6.66 3.24 2.75 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.63 0.575 2.63 0.575 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 14.025 3.62 14.025 2.63 14.255 2.63 14.255 3.62 14.42 3.62 15.12 3.62 15.12 4.22 14.42 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.18 0.865 6.38 0.865 6.38 0.53 14.42 0.53 14.42 0.76 6.61 0.76 6.61 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_2
