# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.56 1.79 3.87 1.79 3.87 2.12 1.56 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.16 1.145 1.16 1.145 2.35 4.12 2.35 4.12 1.79 4.9 1.79 4.9 2.12 4.38 2.12 4.38 2.68 0.825 2.68  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.72 1.19 6.485 1.19 6.485 1.325 8.38 1.325 8.38 1.19 9.42 1.19 9.42 2.19 8.865 2.19 8.865 1.555 6.04 1.555 6.04 2.15 5.72 2.15  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.28 1.8 8.32 1.8 8.32 2.14 6.28 2.14  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.8374 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.13 2.92 4.63 2.92 4.63 2.37 5.15 2.37 5.15 1.56 1.53 1.56 1.53 0.99 1.87 0.99 1.87 1.22 3.77 1.22 3.77 0.99 4.11 0.99 4.11 1.22 5.48 1.22 5.48 2.38 8.56 2.38 8.56 3.275 8.33 3.275 8.33 2.68 6.52 2.68 6.52 3.275 6.29 3.275 6.29 2.68 4.86 2.68 4.86 3.28 2.13 3.28  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.485 0.575 2.485 0.575 3.62 5.115 3.62 5.115 3.205 5.455 3.205 5.455 3.62 7.255 3.62 7.255 3.205 7.595 3.205 7.595 3.62 9.35 3.62 9.35 2.595 9.58 2.595 9.58 3.62 9.645 3.62 10.08 3.62 10.08 4.22 9.645 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 7.595 0.3 7.595 0.635 7.255 0.635 7.255 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.53 6.965 0.53 6.965 0.865 7.85 0.865 7.85 0.53 9.645 0.53 9.645 0.76 8.08 0.76 8.08 1.095 6.735 1.095 6.735 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_2
