* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
M_tn0 VSS E net4 VPW nmos_5p0 W=4.6e-07 L=6e-07
M_tn8 net7 net4 VSS VPW nmos_5p0 W=3.9e-07 L=6e-07
M_tn4 VSS D net3 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn5 net5 net7 net3 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn1 net2 net4 net5 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn2 net2 net6 VSS VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn3 net6 net5 VSS VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn6 Q net5 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_tp0 VDD E net4 VNW pmos_5p0 W=9.2e-07 L=5e-07
M_tp8 net7 net4 VDD VNW pmos_5p0 W=6.25e-07 L=5e-07
M_tp5 VDD D net1 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp4 net1 net4 net5 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp2 net5 net7 net0 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp1 net0 net6 VDD VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp3 net6 net5 VDD VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp6 Q net5 VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
