* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
M_i_4_1 VSS A3 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_1 net_0 A2 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2_1 VSS A1 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 A1 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_0 VSS A2 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_4_0 net_0 A3 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_0 ZN B2 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 B1 ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_1 ZN B1 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 B2 ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_9_1 net_3_0 A3 VDD VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_8_1 net_2_0 A2 net_3_0 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_7_1 ZN A1 net_2_0 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_7_0 net_2_1 A1 ZN VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_8_0 net_3_1 A2 net_2_1 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_9_0 VDD A3 net_3_1 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_6_0 net_1_0 B2 VDD VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_5_0 ZN B1 net_1_0 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_5_1 net_1_1 B1 ZN VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_6_1 VDD B2 net_1_1 VNW pmos_5p0 W=1.095e-06 L=5e-07
.ENDS
