# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.84 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.625 1.77 1.625 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.785 7.72 1.785 7.72 2.15 4.57 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.2676 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.505 2.53 16.325 2.53 16.85 2.53 16.85 1.155 15.74 1.155 15.74 1.135 13.51 1.135 13.51 0.63 13.74 0.63 13.74 0.865 15.75 0.865 15.75 0.635 15.98 0.635 15.98 0.865 17.99 0.865 17.99 0.635 18.22 0.635 18.22 0.865 20.23 0.865 20.23 0.635 20.46 0.635 20.46 1.135 18.315 1.135 18.315 1.155 17.34 1.155 17.34 2.53 19.91 2.53 19.91 3.38 19.68 3.38 19.68 2.83 17.87 2.83 17.87 3.38 17.64 3.38 17.64 2.83 16.325 2.83 15.83 2.83 15.83 3.38 15.6 3.38 15.6 2.83 13.745 2.83 13.745 3.38 13.505 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.535 3.62 1.535 3.285 1.88 3.285 1.88 3.62 4.955 3.62 4.955 3.445 5.295 3.445 5.295 3.62 7.555 3.62 7.555 3.445 7.915 3.445 7.915 3.62 10.1 3.62 10.1 2.665 10.33 2.665 10.33 3.62 12.34 3.62 12.34 2.665 12.57 2.665 12.57 3.62 14.58 3.62 14.58 3.23 14.81 3.23 14.81 3.62 16.325 3.62 16.62 3.62 16.62 3.23 16.85 3.23 16.85 3.62 18.66 3.62 18.66 3.23 18.89 3.23 18.89 3.62 20.46 3.62 20.7 3.62 20.7 2.53 20.93 2.53 20.93 3.62 21.14 3.62 21.84 3.62 21.84 4.22 21.14 4.22 20.46 4.22 16.325 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.84 -0.3 21.84 0.3 21.58 0.3 21.58 1.015 21.35 1.015 21.35 0.3 19.395 0.3 19.395 0.635 19.055 0.635 19.055 0.3 17.155 0.3 17.155 0.635 16.815 0.635 16.815 0.3 14.915 0.3 14.915 0.635 14.575 0.635 14.575 0.3 12.62 0.3 12.62 0.865 12.39 0.865 12.39 0.3 10.38 0.3 10.38 0.865 10.15 0.865 10.15 0.3 8.195 0.3 8.195 0.635 7.855 0.635 7.855 0.3 5.295 0.3 5.295 0.53 5.01 0.53 5.01 0.3 1.61 0.3 1.61 0.76 1.38 0.76 1.38 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.575 2.57 1.955 2.57 1.955 1.225 0.26 1.225 0.26 0.675 0.49 0.675 0.49 0.99 2.185 0.99 2.185 2.09 3.345 2.09 3.345 2.32 2.185 2.32 2.185 2.8 0.805 2.8 0.805 3.38 0.575 3.38  ;
        POLYGON 6.105 2.525 8.5 2.525 8.5 1.555 6.515 1.555 6.515 0.99 6.935 0.99 6.935 1.325 8.73 1.325 8.73 1.625 12.145 1.625 12.145 1.955 8.73 1.955 8.73 2.755 6.58 2.755 6.58 2.78 6.105 2.78  ;
        POLYGON 2.5 0.53 4.78 0.53 4.78 0.76 5.77 0.76 5.77 0.53 7.395 0.53 7.395 0.865 9.03 0.865 9.03 0.53 9.26 0.53 9.26 0.865 9.635 0.865 9.635 1.095 11.27 1.095 11.27 0.53 11.5 0.53 11.5 1.095 12.62 1.095 12.62 1.365 15.48 1.365 15.48 1.595 12.39 1.595 12.39 1.325 9.405 1.325 9.405 1.095 7.165 1.095 7.165 0.76 6 0.76 6 0.99 4.55 0.99 4.55 0.76 3.22 0.76 3.22 1.575 3.865 1.575 3.865 2.89 3.635 2.89 3.635 1.805 2.99 1.805 2.99 0.885 2.5 0.885  ;
        POLYGON 2.52 3.125 4.095 3.125 4.095 1.345 3.775 1.345 3.775 0.99 4.135 0.99 4.135 1.115 4.325 1.115 4.325 2.985 5.875 2.985 5.875 3.055 6.81 3.055 6.81 2.985 9.025 2.985 9.025 2.185 12.39 2.185 12.39 1.96 16.325 1.96 16.325 2.195 12.62 2.195 12.62 2.415 11.45 2.415 11.45 3.26 11.22 3.26 11.22 2.415 9.365 2.415 9.365 3.215 7.325 3.215 7.325 3.355 5.525 3.355 5.525 3.215 4.725 3.215 4.725 3.355 2.52 3.355  ;
        POLYGON 18.165 1.96 20.46 1.96 20.46 2.195 18.165 2.195  ;
        POLYGON 18.505 1.365 21.14 1.365 21.14 1.595 18.505 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_8
