# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 7.184 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.765 3.79 1.765 3.79 2.15 0.63 2.15  ;
        POLYGON 5.33 1.765 8.96 1.765 8.96 2.15 5.33 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.41 4.57 2.41 4.57 1.535 1.365 1.535 1.365 0.7 1.595 0.7 1.595 1.215 3.605 1.215 3.605 0.7 3.835 0.7 3.835 1.215 5.845 1.215 5.845 0.7 6.075 0.7 6.075 1.215 8.085 1.215 8.085 0.7 8.315 0.7 8.315 1.535 4.95 1.535 4.95 2.41 8.215 2.41 8.215 3.38 7.985 3.38 7.985 2.725 5.975 2.725 5.975 3.38 5.745 3.38 5.745 2.725 3.735 2.725 3.735 3.38 3.505 3.38 3.505 2.73 1.495 2.73 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.55 0.475 2.55 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 4.57 3.62 4.57 2.965 4.91 2.965 4.91 3.62 6.81 3.62 6.81 2.965 7.15 2.965 7.15 3.62 9.105 3.62 9.105 2.55 9.335 2.55 9.335 3.62 10.08 3.62 10.08 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.435 0.3 9.435 1.04 9.205 1.04 9.205 0.3 7.25 0.3 7.25 0.985 6.91 0.985 6.91 0.3 5.01 0.3 5.01 0.985 4.67 0.985 4.67 0.3 2.77 0.3 2.77 0.985 2.43 0.985 2.43 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_8
