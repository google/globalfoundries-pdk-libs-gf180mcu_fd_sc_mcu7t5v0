# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 0.55 3.24 0.55 3.24 2.15 2.92 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 0.55 3.8 0.55 3.8 1.8 4.545 1.8 4.545 2.15 3.48 2.15  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.55 2.12 0.55 2.12 2.15 1.8 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.085 1.005 1.085 1.005 1.77 1.57 1.77 1.57 2.15 0.61 2.15  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 0.585 2.68 0.585 2.68 2.38 3.89 2.38 3.89 2.71 2.35 2.71  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.33 3.62 1.33 3.04 1.56 3.04 1.56 3.62 4.675 3.62 5.04 3.62 5.04 4.22 4.675 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.62 0.3 4.62 0.905 4.39 0.905 4.39 0.3 0.54 0.3 0.54 0.725 0.31 0.725 0.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.255 2.53 2.05 2.53 2.05 3.145 4.335 3.145 4.335 2.53 4.675 2.53 4.675 3.38 1.82 3.38 1.82 2.76 0.595 2.76 0.595 3.38 0.255 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_1
