* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 D RN SETN CLK Q VDD VNW VPW VSS
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp10 net3 cki net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS
