* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_14 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_15 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_18 I3 I2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_19 VSS A3 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_10 Z_neg I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 net_2 A3 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 VSS I2 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_1 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_0 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_16 net_4 A2 I VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_17 VDD A1 net_4 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_20 net_5 I2 I3 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_21 VDD A3 net_5 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_13 net_3 I3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11 Z_neg A3 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_12 net_3 I2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS
