# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.54 1.02 1.54 1.02 2.81 0.66 2.81  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.54 2.14 1.54 2.14 3.37 1.78 3.37  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 0.555 3.87 0.555 3.87 3.38 3.45 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.225 0.475 3.225 0.475 3.62 2.605 3.62 2.605 2.53 2.835 2.53 2.835 3.62 3.175 3.62 4.48 3.62 4.48 4.22 3.175 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.735 0.3 2.735 0.765 2.505 0.765 2.505 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.805 0.475 0.805 0.475 1.055 3.175 1.055 3.175 1.985 2.945 1.985 2.945 1.29 1.495 1.29 1.495 3.325 1.265 3.325 1.265 1.29 0.245 1.29  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_1
