# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.64 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.095 1.77 6.785 1.77 6.785 2.15 5.095 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 19.65 1.77 19.65 2.16 17.45 2.16  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.734 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.33 1.625 11.86 1.625 12.325 1.625 12.325 0.65 12.755 0.65 12.755 1.625 16.615 1.625 17.11 1.625 17.11 1.855 16.615 1.855 11.86 1.855 7.33 1.855  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5972 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.79 1.92 22.785 1.92 23.03 1.92 23.03 1.135 20.805 1.135 20.805 0.53 21.035 0.53 21.035 0.905 23.03 0.905 23.03 0.53 23.41 0.53 23.41 3.37 23.03 3.37 23.03 2.24 22.785 2.24 21.26 2.24 21.26 3.37 20.79 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.675 1.92 3.915 1.92 3.915 3.37 3.46 3.37 3.46 2.24 1.675 2.24 1.675 3.37 1.215 3.37 1.215 0.53 1.675 0.53 1.675 0.905 3.685 0.905 3.685 0.53 3.915 0.53 3.915 1.135 1.675 1.135  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.325 3.62 0.325 2.65 0.555 2.65 0.555 3.62 2.565 3.62 2.565 2.65 2.795 2.65 2.795 3.62 4.805 3.62 4.805 3.16 5.035 3.16 5.035 3.62 8.11 3.62 10.23 3.62 10.23 3.005 10.57 3.005 10.57 3.62 11.93 3.62 12.765 3.62 12.765 2.67 12.995 2.67 12.995 3.62 14.99 3.62 14.99 3.005 15.33 3.005 15.33 3.62 16.57 3.62 19.585 3.62 19.585 3.16 19.815 3.16 19.815 3.62 21.925 3.62 21.925 2.56 22.155 2.56 22.155 3.62 22.785 3.62 24.165 3.62 24.165 2.56 24.395 2.56 24.395 3.62 24.64 3.62 24.64 4.22 22.785 4.22 16.57 4.22 11.93 4.22 8.11 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.64 -0.3 24.64 0.3 24.395 0.3 24.395 0.765 24.165 0.765 24.165 0.3 22.21 0.3 22.21 0.67 21.87 0.67 21.87 0.3 19.915 0.3 19.915 0.765 19.685 0.765 19.685 0.3 15.33 0.3 15.33 0.915 14.99 0.915 14.99 0.3 13.215 0.3 13.215 1.135 12.985 1.135 12.985 0.3 10.57 0.3 10.57 0.915 10.23 0.915 10.23 0.3 5.09 0.3 5.09 0.675 4.75 0.675 4.75 0.3 2.85 0.3 2.85 0.675 2.505 0.675 2.505 0.3 0.555 0.3 0.555 0.87 0.325 0.87 0.325 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.79 2.545 8.11 2.545 8.11 2.775 4.56 2.775 4.56 1.67 1.915 1.67 1.915 1.44 4.56 1.44 4.56 0.905 7.77 0.905 7.77 0.78 8.11 0.78 8.11 1.14 4.79 1.14  ;
        POLYGON 8.945 0.795 9.175 0.795 9.175 1.145 11.63 1.145 11.63 0.795 11.86 0.795 11.86 1.375 8.945 1.375  ;
        POLYGON 8.99 2.545 11.93 2.545 11.93 2.83 11.59 2.83 11.59 2.775 9.33 2.775 9.33 2.83 8.99 2.83  ;
        POLYGON 13.74 2.545 16.57 2.545 16.57 2.775 13.74 2.775  ;
        POLYGON 13.705 0.81 13.935 0.81 13.935 1.145 16.385 1.145 16.385 0.81 16.615 0.81 16.615 1.375 13.705 1.375  ;
        POLYGON 8.38 2.085 17.165 2.085 17.165 2.55 20.125 2.55 20.125 1.365 17.505 1.365 17.505 0.81 17.735 0.81 17.735 1.135 20.355 1.135 20.355 1.44 22.785 1.44 22.785 1.67 20.355 1.67 20.355 2.785 16.935 2.785 16.935 2.315 8.38 2.315  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_4
