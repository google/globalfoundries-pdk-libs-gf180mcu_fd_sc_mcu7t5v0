* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1_1 net_0_0 A2 VSS VPW nmos_5p0 W=7.8e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=7.8e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=7.8e-07 L=6e-07
M_i_1_0 VSS A2 net_0_1 VPW nmos_5p0 W=7.8e-07 L=6e-07
M_i_2_0 ZN B VSS VPW nmos_5p0 W=5.15e-07 L=6e-07
M_i_3_0 VSS C ZN VPW nmos_5p0 W=5.15e-07 L=6e-07
M_i_3_1 ZN C VSS VPW nmos_5p0 W=5.15e-07 L=6e-07
M_i_2_1 VSS B ZN VPW nmos_5p0 W=5.15e-07 L=6e-07
M_i_5_1 ZN A2 net_1 VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_4_1 net_1 A1 ZN VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_4_0 ZN A1 net_1 VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_5_0 net_1 A2 ZN VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_6_0 net_2_0 B net_1 VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_7_0 VDD C net_2_0 VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_7_1 net_2_1 C VDD VNW pmos_5p0 W=1.14e-06 L=5e-07
M_i_6_1 net_1 B net_2_1 VNW pmos_5p0 W=1.14e-06 L=5e-07
.ENDS
