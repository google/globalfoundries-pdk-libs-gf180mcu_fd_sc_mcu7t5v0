# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0995 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.775 1.77 2.34 1.77 2.34 1.16 2.68 1.16 2.68 2.15 1.775 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0995 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.115 1.77 0.66 1.77 0.66 1.16 1.01 1.16 1.01 2.15 0.115 2.15  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9135 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.91 1.77 3.475 1.77 3.475 1.16 3.815 1.16 3.815 2.15 2.91 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1456 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.24 0.55 2.58 0.55 2.58 0.87 1.545 0.87 1.545 2.725 1.24 2.725  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.57 3.62 3.525 3.62 3.525 2.69 3.755 2.69 3.755 3.62 4.48 3.62 4.48 4.22 2.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 3.855 0.3 3.855 0.765 3.625 0.765 3.625 0.3 0.475 0.3 0.475 0.765 0.245 0.765 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 2.495 0.53 2.495 0.53 3.16 2.23 3.16 2.23 2.495 2.57 2.495 2.57 3.39 0.19 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_1
