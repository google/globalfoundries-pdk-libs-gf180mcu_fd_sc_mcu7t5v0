# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.3 1.06 7.72 1.06 7.72 1.77 8.2 1.77 8.27 1.77 8.27 2.15 8.2 2.15 7.3 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.72 1.06 6.04 1.06 6.04 1.77 6.61 1.77 6.61 2.15 5.72 2.15  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.37 1.77 4.36 1.77 4.36 2.15 2.69 2.15 2.69 3.32 2.37 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.59 1.77 4.61 1.77 5.16 1.77 5.16 1.06 5.48 1.06 5.48 2.15 4.61 2.15 4.59 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.78 1.52 2.14 1.52 2.14 3.32 1.78 3.32  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.66 1.16 1.02 1.16 1.02 2.71 0.66 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5684 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.055 2.9 4.61 2.9 4.755 2.9 4.755 2.74 6.84 2.74 6.84 1.22 6.51 1.22 6.51 0.99 7.07 0.99 7.07 2.74 8.1 2.74 8.1 3.26 6.035 3.26 6.035 2.97 5.065 2.97 5.065 3.26 4.61 3.26 3.055 3.26  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.95 0.575 2.95 0.575 3.62 4.61 3.62 5.445 3.62 5.445 3.2 5.675 3.2 5.675 3.62 8.2 3.62 8.4 3.62 8.4 4.22 8.2 4.22 4.61 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 2.715 0.3 2.715 0.76 2.485 0.76 2.485 0.3 0.475 0.3 0.475 0.76 0.245 0.76 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 0.53 1.595 0.53 1.595 0.99 4.61 0.99 4.61 1.22 1.365 1.22  ;
        POLYGON 3.15 0.53 8.2 0.53 8.2 0.76 3.15 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_1
