# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.61 1.015 0.61 1.015 1.625 1.65 1.625 1.65 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.675 2.21 3.24 2.21 3.48 2.21 3.48 1.3 2.675 1.3 2.675 0.57 2.905 0.57 2.905 1.065 3.8 1.065 3.8 2.7 3.24 2.7 2.905 2.7 2.905 3.39 2.675 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.405 3.62 1.405 3.01 1.745 3.01 1.745 3.62 3.24 3.62 3.64 3.62 3.64 3.01 3.98 3.01 3.98 3.62 4.48 3.62 4.48 4.22 3.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 4.08 0.3 4.08 0.765 3.74 0.765 3.74 0.3 1.745 0.3 1.745 0.765 1.405 0.765 1.405 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.57 0.475 0.57 0.475 2.39 1.9 2.39 1.9 1.55 3.24 1.55 3.24 1.89 2.13 1.89 2.13 2.625 0.475 2.625 0.475 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_2
