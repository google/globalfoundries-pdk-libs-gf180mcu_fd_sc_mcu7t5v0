# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.485 1.78 16.51 1.78 18.175 1.78 18.175 2.12 16.51 2.12 16.485 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.835 1.78 13.735 1.78 13.735 2.13 11.835 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.97 1.01 0.97 1.01 2.95 0.705 2.95  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.505 0.55 4.935 0.55 4.935 1.8 5.755 1.8 5.755 2.15 4.505 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.255 1.8 3.3 1.8 3.3 1.24 3.7 1.24 3.7 2.25 2.255 2.25  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.17 1.305 9.535 1.305 9.535 1.77 9.95 1.77 10.535 1.77 10.535 3.32 10.165 3.32 10.165 2.15 9.95 2.15 9.17 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.7592 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 0.6 6.6 0.6 6.6 2.855 6.23 2.855  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.575 0.475 2.575 0.475 3.62 1.65 3.62 5.01 3.62 5.01 2.845 5.35 2.845 5.35 3.62 7.405 3.62 7.405 2.57 7.635 2.57 7.635 3.62 8.48 3.62 9.95 3.62 12.905 3.62 12.905 2.845 13.25 2.845 13.25 3.62 15.335 3.62 17.19 3.62 17.19 2.815 17.53 2.815 17.53 3.62 18.695 3.62 19.04 3.62 19.04 4.22 18.695 4.22 15.335 4.22 9.95 4.22 8.48 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 17.575 0.3 17.575 1.145 17.345 1.145 17.345 0.3 13.095 0.3 13.095 1.145 12.865 1.145 12.865 0.3 7.635 0.3 7.635 1.16 7.405 1.16 7.405 0.3 5.395 0.3 5.395 1.16 5.165 1.16 5.165 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 2.95 1.26 2.95  ;
        POLYGON 3.93 0.78 4.275 0.78 4.275 2.87 3.93 2.87  ;
        POLYGON 8.095 2.665 8.48 2.665 8.48 3.005 7.865 3.005 7.865 2.275 7.095 2.275 7.095 3.39 5.67 3.39 5.67 2.615 4.735 2.615 4.735 3.33 2.71 3.33 2.71 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.91 0.845 2.91 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 3.05 2.74 3.05 3.1 4.505 3.1 4.505 2.38 5.9 2.38 5.9 3.155 6.865 3.155 6.865 2.045 7.865 2.045 7.865 0.79 8.48 0.79 8.48 1.13 8.095 1.13  ;
        POLYGON 8.325 1.46 8.71 1.46 8.71 0.845 9.95 0.845 9.95 1.075 8.94 1.075 8.94 2.72 9.88 2.72 9.88 2.95 8.71 2.95 8.71 1.82 8.325 1.82  ;
        POLYGON 11.595 2.575 12.075 2.575 12.075 2.925 11.345 2.925 11.345 0.795 12.075 0.795 12.075 1.145 11.595 1.145  ;
        POLYGON 13.985 0.78 14.215 0.78 14.215 2.925 13.985 2.925  ;
        POLYGON 10.885 0.78 11.115 0.78 11.115 3.16 12.36 3.16 12.36 2.38 13.73 2.38 13.73 3.16 15.005 3.16 15.005 0.78 15.335 0.78 15.335 3.39 13.5 3.39 13.5 2.615 12.59 2.615 12.59 3.39 10.885 3.39  ;
        POLYGON 15.565 0.85 16.51 0.85 16.51 1.08 15.795 1.08 15.795 2.815 16.425 2.815 16.425 3.045 15.565 3.045  ;
        POLYGON 16.025 1.675 16.255 1.675 16.255 2.355 18.465 2.355 18.465 0.78 18.695 0.78 18.695 3.14 18.36 3.14 18.36 2.585 16.025 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_2
