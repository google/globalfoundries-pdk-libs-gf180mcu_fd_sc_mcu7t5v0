# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.65 1.715 3.51 1.715 3.51 2.15 0.65 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.7312 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.845 2.33 8.27 2.33 8.84 2.33 8.84 1.42 5.845 1.42 5.845 0.675 6.105 0.675 6.105 1.04 8.085 1.04 8.085 0.675 8.315 0.675 8.315 1.04 10.325 1.04 10.325 0.675 10.555 0.675 10.555 1.04 12.565 1.04 12.565 0.675 12.795 0.675 12.795 1.42 9.64 1.42 9.64 2.33 12.695 2.33 12.695 3.38 12.465 3.38 12.465 2.71 10.455 2.71 10.455 3.38 10.225 3.38 10.225 2.71 8.27 2.71 8.215 2.71 8.215 3.38 7.985 3.38 7.985 2.71 6.075 2.71 6.075 3.38 5.845 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.385 3.62 2.385 3.04 2.615 3.04 2.615 3.62 4.625 3.62 4.625 2.57 4.855 2.57 4.855 3.62 6.865 3.62 6.865 3.04 7.095 3.04 7.095 3.62 8.27 3.62 9.105 3.62 9.105 3.04 9.335 3.04 9.335 3.62 11.345 3.62 11.345 3.04 11.575 3.04 11.575 3.62 13.54 3.62 13.585 3.62 13.585 2.57 13.815 2.57 13.815 3.62 14.56 3.62 14.56 4.22 13.54 4.22 8.27 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.97 0.3 13.97 0.765 13.63 0.765 13.63 0.3 11.73 0.3 11.73 0.765 11.39 0.765 11.39 0.3 9.49 0.3 9.49 0.765 9.15 0.765 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 3.98 2.53 3.98 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 4.315 1.015 4.315 1.685 8.27 1.685 8.27 2.025 4.315 2.025 4.315 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 10.34 1.685 13.54 1.685 13.54 2.03 10.34 2.03  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_8
