# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 1.77 4.69 1.77 4.69 1.45 12.42 1.45 12.42 1.68 4.92 1.68 4.92 2.15 3.48 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 2.22 5.42 2.22 5.42 1.91 5.92 1.91 5.92 2.22 8.86 2.22 8.86 1.91 10.22 1.91 10.22 2.22 12.97 2.22 12.97 1.725 13.89 1.725 13.89 2.45 6.775 2.45 6.775 2.71 5.15 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.68 3.24 1.68 3.24 2.15 0.62 2.15  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.89 1.785 19.15 1.785 19.15 2.12 14.89 2.12  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.0289 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.13 2.7 14.12 2.7 14.12 1.22 1.31 1.22 1.31 0.99 14.44 0.99 14.44 2.36 18.43 2.36 18.43 2.93 7.13 2.93  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.53 3.62 1.53 3.285 1.87 3.285 1.87 3.62 3.77 3.62 3.77 3.285 4.11 3.285 4.11 3.62 14.1 3.62 14.47 3.62 14.47 3.285 14.81 3.285 14.81 3.62 16.61 3.62 16.61 3.285 16.95 3.285 16.95 3.62 18.855 3.62 18.855 2.57 19.085 2.57 19.085 3.62 19.2 3.62 19.6 3.62 19.6 4.22 19.2 4.22 14.1 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.6 -0.3 19.6 0.3 18.07 0.3 18.07 0.635 17.73 0.635 17.73 0.3 15.83 0.3 15.83 0.635 15.49 0.635 15.49 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.57 4.59 2.57 4.59 3.16 14.1 3.16 14.1 3.39 4.36 3.39 4.36 2.8 2.935 2.8 2.935 3.38 2.705 3.38 2.705 2.8 0.575 2.8 0.575 3.38 0.345 3.38  ;
        POLYGON 0.18 0.53 15.21 0.53 15.21 0.865 19.2 0.865 19.2 1.095 14.98 1.095 14.98 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_4
