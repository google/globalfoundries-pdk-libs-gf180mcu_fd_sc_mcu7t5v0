# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 1.765 4.39 1.765 4.39 2.19 3.095 2.19  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.315 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.155 1.21 20.035 1.21 20.035 0.665 20.7 0.665 20.7 1.02 20.41 1.02 20.41 1.635 19.155 1.635  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.11375 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.46 0.6 23.98 0.6 23.98 3.36 23.46 3.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 10.125 3.62 10.62 3.62 13.12 3.62 13.12 3 13.46 3 13.46 3.62 14.645 3.62 15.135 3.62 15.135 2.665 15.365 2.665 15.365 3.62 16.385 3.62 19.48 3.62 19.48 2.845 19.82 2.845 19.82 3.62 21.345 3.62 21.675 3.62 21.675 2.57 21.905 2.57 21.905 3.62 22.445 3.62 22.445 2.56 22.675 2.56 22.675 3.62 23.145 3.62 24.535 3.62 24.535 2.56 24.765 2.56 24.765 3.62 25.2 3.62 25.2 4.22 23.145 4.22 21.345 4.22 16.385 4.22 14.645 4.22 10.62 4.22 10.125 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 24.865 0.3 24.865 0.925 24.635 0.925 24.635 0.3 22.625 0.3 22.625 0.925 22.395 0.925 22.395 0.3 19.7 0.3 19.7 0.915 19.36 0.915 19.36 0.3 14.71 0.3 14.71 0.915 14.37 0.915 14.37 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 4.845 2.745 4.845 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.895 3.16 9.895 2.645 10.125 2.645 10.125 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 5.075 2.655 5.075 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.375 1.26 6.375 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.97 9.925 0.97 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.605 0.76 6.605 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.62 1.8 10.62 2.035 9.115 2.035 9.115 2.845 8.885 2.845  ;
        POLYGON 11.935 2.53 14.645 2.53 14.645 3.005 14.415 3.005 14.415 2.76 12.165 2.76 12.165 3.005 11.935 3.005  ;
        POLYGON 10.915 2.065 11.045 2.065 11.045 0.63 11.275 0.63 11.275 2.065 11.965 2.065 11.965 1.61 15.37 1.61 15.37 1.84 12.195 1.84 12.195 2.295 11.145 2.295 11.145 3.125 10.915 3.125  ;
        POLYGON 12.46 2.07 15.71 2.07 15.71 0.99 16.05 0.99 16.05 2.07 16.385 2.07 16.385 3.035 16.155 3.035 16.155 2.3 12.46 2.3  ;
        POLYGON 11.505 1.145 14.98 1.145 14.98 0.53 17.845 0.53 17.845 2.06 17.99 2.06 17.99 2.4 17.615 2.4 17.615 0.76 16.6 0.76 16.6 1.735 16.37 1.735 16.37 0.76 15.21 0.76 15.21 1.375 11.735 1.375 11.735 1.72 11.505 1.72  ;
        POLYGON 18.075 0.79 18.305 0.79 18.305 1.51 18.45 1.51 18.45 2.42 18.57 2.42 18.57 2.93 18.22 2.93 18.22 1.745 18.075 1.745  ;
        POLYGON 16.83 0.99 17.385 0.99 17.385 2.69 17.46 2.69 17.46 3.16 18.845 3.16 18.845 2.385 20.425 2.385 20.425 3.155 21.115 3.155 21.115 2.03 21.345 2.03 21.345 3.39 20.195 3.39 20.195 2.615 19.075 2.615 19.075 3.39 17.155 3.39 17.155 1.22 16.83 1.22  ;
        POLYGON 18.68 1.68 18.91 1.68 18.91 1.925 20.655 1.925 20.655 1.405 21.675 1.405 21.675 0.81 21.905 0.81 21.905 1.405 23.145 1.405 23.145 2.25 22.915 2.25 22.915 1.635 20.885 1.635 20.885 2.86 20.655 2.86 20.655 2.155 18.68 2.155  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
