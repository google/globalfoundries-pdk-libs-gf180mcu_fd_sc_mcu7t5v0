# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.835 1.465 8.47 1.465 8.47 1.24 9.63 1.24 9.63 1.56 8.745 1.56 8.745 1.695 6.835 1.695  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.69 1.75 6.605 1.75 6.605 1.93 8.975 1.93 8.975 1.8 9.63 1.8 9.63 2.16 5.69 2.16  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 1.825 1.275 1.825 1.275 1.93 3.45 1.93 3.45 1.825 4.615 1.825 4.615 2.16 0.385 2.16  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 1.265 1.735 1.265 1.735 1.465 3.22 1.465 3.22 1.695 1.505 1.695 1.505 1.565 0.385 1.565  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.631 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.53 2.205 0.53 2.205 1.005 3.005 1.005 3.005 0.53 4.625 0.53 4.625 1.005 5.425 1.005 5.425 0.53 7.045 0.53 7.045 1.005 7.845 1.005 7.845 0.53 8.95 0.53 8.95 0.975 8.145 0.975 8.145 1.235 6.815 1.235 6.815 0.975 5.655 0.975 5.655 1.235 5.46 1.235 5.46 2.39 7.79 2.39 7.79 2.665 5.13 2.665 5.13 1.235 4.395 1.235 4.395 0.975 3.235 0.975 3.235 1.235 1.975 1.235 1.975 0.975 1.17 0.975  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.44 3.62 2.44 2.935 2.67 2.935 2.67 3.62 9.7 3.62 10.08 3.62 10.08 4.22 9.7 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.855 0.3 9.855 0.775 9.515 0.775 9.515 0.3 7.615 0.3 7.615 0.775 7.275 0.775 7.275 0.3 5.195 0.3 5.195 0.775 4.855 0.775 4.855 0.3 2.775 0.3 2.775 0.775 2.435 0.775 2.435 0.3 0.535 0.3 0.535 0.775 0.195 0.775 0.195 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.35 2.39 4.615 2.39 4.615 2.965 9.47 2.965 9.47 2.53 9.7 2.53 9.7 3.38 9.47 3.38 9.47 3.195 4.385 3.195 4.385 2.625 0.58 2.625 0.58 3.38 0.35 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor4_2
