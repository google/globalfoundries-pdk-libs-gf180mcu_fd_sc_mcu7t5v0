# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.85 1.8 4.39 1.8 4.39 2.12 2.85 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 1.77 2.35 1.77 2.35 1.325 4.85 1.325 4.85 1.77 6.07 1.77 6.07 2.12 4.62 2.12 4.62 1.555 2.6 1.555 2.6 2.135 1.535 2.135  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.56 1.145 1.56 1.145 2.365 6.3 2.365 6.3 1.56 6.6 1.56 6.6 2.595 6.16 2.595 6.16 2.68 0.825 2.68  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.45 1.8 10.59 1.8 10.59 2.12 8.45 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.56 1.785 7.88 1.785 7.88 2.365 11.215 2.365 11.215 1.56 11.535 1.56 11.535 2.68 8.12 2.68 8.12 2.595 7.56 2.595  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3774 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 2.92 6.41 2.92 6.41 2.825 6.84 2.825 6.84 0.99 10.84 0.99 10.84 1.22 7.16 1.22 7.16 2.825 7.75 2.825 7.75 2.92 10.17 2.92 10.17 3.24 7.5 3.24 7.5 3.055 6.66 3.055 6.66 3.24 3.365 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.65 0.575 2.65 0.575 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 11.785 3.62 11.785 2.65 12.015 2.65 12.015 3.62 12.18 3.62 12.88 3.62 12.88 4.22 12.18 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 6.37 0.865 6.37 0.53 12.18 0.53 12.18 0.76 6.6 0.76 6.6 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_2
