* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
M_i_8 net_2 A2 I VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_9 VSS A1 net_2 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_4 net_0 I VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_2 Z_neg A1 net_0 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3 net_0 A2 Z_neg VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_10 I A2 VDD VNW pmos_5p0 W=3.85e-07 L=5e-07
M_i_11 VDD A1 I VNW pmos_5p0 W=3.85e-07 L=5e-07
M_i_7 Z_neg I VDD VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_5 net_1 A1 Z_neg VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_6 VDD A2 net_1 VNW pmos_5p0 W=1.095e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
