# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5305 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1565 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.56 1.22 15.59 1.22 15.59 1.67 14.56 1.67  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.794 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.61 2.09 19.93 2.09 20.26 2.09 20.26 1.29 19.665 1.29 19.665 0.55 20.06 0.55 20.06 1.06 20.62 1.06 20.62 2.32 20.06 2.32 20.06 3.38 19.93 3.38 19.61 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.155 3.62 3.05 3.62 3.05 3.005 3.39 3.005 3.39 3.62 7.29 3.62 7.29 3.24 7.63 3.24 7.63 3.62 9.825 3.62 9.825 2.885 10.055 2.885 10.055 3.62 11.67 3.62 14.11 3.62 14.11 2.945 14.45 2.945 14.45 3.62 16.745 3.62 16.745 2.6 16.975 2.6 16.975 3.62 17.47 3.62 18.645 3.62 18.645 2.57 18.875 2.57 18.875 3.62 19.93 3.62 20.685 3.62 20.685 2.57 20.915 2.57 20.915 3.62 21.28 3.62 21.28 4.22 19.93 4.22 17.47 4.22 11.67 4.22 2.155 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 21.015 0.3 21.015 0.765 20.785 0.765 20.785 0.3 18.775 0.3 18.775 0.765 18.545 0.765 18.545 0.3 16.99 0.3 16.99 1.08 16.65 1.08 16.65 0.3 7.81 0.3 7.81 1.09 7.47 1.09 7.47 0.3 3.455 0.3 3.455 1.145 3.225 1.145 3.225 0.3 1.65 0.3 1.65 0.935 1.31 0.935 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.36 1.925 2.36 1.925 1.395 0.245 1.395 0.245 0.66 0.475 0.66 0.475 1.165 2.155 1.165 2.155 2.595 0.575 2.595 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 2.52 4.86 2.52 4.86 1.095 4.29 1.095 4.29 0.865 5.09 0.865 5.09 2.75 4.29 2.75  ;
        POLYGON 5.365 0.865 5.85 0.865 5.85 1.395 8.29 1.395 8.29 1.63 5.595 1.63 5.595 2.71 5.365 2.71  ;
        POLYGON 6.63 1.965 9.825 1.965 9.825 0.81 10.055 0.81 10.055 1.93 11.23 1.93 11.23 2.655 10.89 2.655 10.89 2.195 8.87 2.195 8.87 2.655 8.53 2.655 8.53 2.195 6.63 2.195  ;
        POLYGON 2.385 0.66 2.715 0.66 2.715 2.545 3.85 2.545 3.85 3.12 5.94 3.12 5.94 2.65 8.205 2.65 8.205 2.885 9.1 2.885 9.1 2.425 10.515 2.425 10.515 3.065 11.67 3.065 11.67 3.295 10.285 3.295 10.285 2.655 9.33 2.655 9.33 3.115 7.975 3.115 7.975 2.88 6.23 2.88 6.23 3.36 3.62 3.36 3.62 2.775 2.715 2.775 2.715 3.3 2.385 3.3  ;
        POLYGON 13.395 1.965 15.73 1.965 15.73 2.655 15.38 2.655 15.38 2.195 13.395 2.195 13.395 2.71 13.165 2.71 13.165 1.075 12.01 1.075 12.01 0.795 14.295 0.795 14.295 1.135 13.395 1.135  ;
        POLYGON 10.945 0.81 11.175 0.81 11.175 1.355 12.375 1.355 12.375 2.94 13.625 2.94 13.625 2.48 14.985 2.48 14.985 2.885 16.15 2.885 16.15 1.96 17.47 1.96 17.47 2.195 16.38 2.195 16.38 3.12 14.755 3.12 14.755 2.715 13.855 2.715 13.855 3.175 12.145 3.175 12.145 1.585 10.945 1.585  ;
        POLYGON 15.99 1.385 17.825 1.385 17.825 0.795 18.055 0.795 18.055 1.605 19.93 1.605 19.93 1.835 17.995 1.835 17.995 2.875 17.765 2.875 17.765 1.615 15.99 1.615  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
