# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.96 1.45 6.79 1.45 6.79 1.77 8.31 1.77 8.31 2.12 6.54 2.12 6.54 1.68 1.96 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.91 6.205 1.91 6.205 2.36 8.54 2.36 8.54 1.77 9.41 1.77 9.41 2.12 8.88 2.12 8.88 2.68 5.955 2.68 5.955 2.14 0.62 2.14  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.2 1.325 12.93 1.325 12.93 1.22 15.08 1.22 15.08 1.325 17.76 1.325 17.76 1.555 10.52 1.555 10.52 2.425 10.2 2.425  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.75 1.8 16.84 1.8 16.84 2.12 10.75 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.279 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.65 2.475 2.99 2.475 2.99 2.92 4.39 2.92 4.39 2.795 5.725 2.795 5.725 2.92 9.09 2.92 9.09 2.795 9.64 2.795 9.64 1.22 1.52 1.22 1.52 0.99 9.96 0.99 9.96 2.795 17.45 2.795 17.45 3.24 16.4 3.24 16.4 3.055 15.56 3.055 15.56 3.24 14.36 3.24 14.36 3.055 13.52 3.055 13.52 3.24 12.32 3.24 12.32 3.055 11.48 3.055 11.48 3.24 10.175 3.24 10.175 3.025 9.34 3.025 9.34 3.24 5.475 3.24 5.475 3.025 4.64 3.025 4.64 3.24 2.99 3.24 2.99 3.325 2.65 3.325  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.89 3.62 4.89 3.285 5.23 3.285 5.23 3.62 9.59 3.62 9.59 3.285 9.93 3.285 9.93 3.62 11.73 3.62 11.73 3.285 12.07 3.285 12.07 3.62 13.77 3.62 13.77 3.285 14.11 3.285 14.11 3.62 15.81 3.62 15.81 3.285 16.15 3.285 16.15 3.62 17.905 3.62 17.905 2.595 18.135 2.595 18.135 3.62 18.2 3.62 18.48 3.62 18.48 4.22 18.2 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.15 0.3 16.15 0.635 15.81 0.635 15.81 0.3 12.07 0.3 12.07 0.635 11.73 0.635 11.73 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.53 10.885 0.53 10.885 0.865 12.32 0.865 12.32 0.53 15.56 0.53 15.56 0.865 18.2 0.865 18.2 1.095 15.33 1.095 15.33 0.76 12.55 0.76 12.55 1.095 10.655 1.095 10.655 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_4
