# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 4.48 3.62 4.48 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.085 2.485 1.085 2.485 0.3 0.475 0.3 0.475 1.085 0.245 1.085 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_8
