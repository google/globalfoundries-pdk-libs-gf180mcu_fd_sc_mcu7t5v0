# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.24 3.16 1.24 3.16 1.56 0.62 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.8 4.03 1.8 4.03 2.12 0.62 2.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6016 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.22 2.36 4.26 2.36 4.26 1.535 3.46 1.535 3.46 1 2.15 1 2.15 0.68 3.82 0.68 3.82 1.265 4.49 1.265 4.49 2.68 3.535 2.68 3.535 3.38 3.305 3.38 3.305 2.68 1.58 2.68 1.58 3.38 1.22 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.285 3.62 2.285 3.085 2.515 3.085 2.515 3.62 4.325 3.62 4.325 3.085 4.555 3.085 4.555 3.62 5.04 3.62 5.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.62 0.3 4.62 0.635 4.26 0.635 4.26 0.3 0.475 0.3 0.475 0.905 0.245 0.905 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_2
