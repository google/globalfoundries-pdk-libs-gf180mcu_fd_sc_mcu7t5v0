# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.405 1.205 4.025 1.205 4.025 1.545 3.405 1.545  ;
        POLYGON 5.645 1.205 6.275 1.205 6.275 1.545 5.645 1.545  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.33 1.78 6.73 1.78 6.73 2.01 3.535 2.01 3.535 2.12 2.33 2.12  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.785 1.575 2.1 1.575 2.1 2.36 3.765 2.36 3.765 2.24 7.41 2.24 7.41 1.665 7.72 1.665 7.72 2.47 3.98 2.47 3.98 2.68 1.785 2.68  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.765 1.21 1.765 1.21 2.92 4.21 2.92 4.21 2.7 7.96 2.7 7.96 1.4 8.885 1.4 8.885 1.63 8.31 1.63 8.31 2.93 4.44 2.93 4.44 3.24 0.87 3.24  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.49 2.36 13.47 2.36 13.73 2.36 13.73 1.56 10.505 1.56 10.505 0.615 10.735 0.615 10.735 1.24 12.745 1.24 12.745 0.615 12.975 0.615 12.975 1.24 13.97 1.24 13.97 2.68 13.47 2.68 12.875 2.68 12.875 3.38 12.645 3.38 12.645 2.68 10.75 2.68 10.75 3.38 10.49 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.555 0.575 2.555 0.575 3.62 9.38 3.62 9.38 2.53 9.61 2.53 9.61 3.62 11.575 3.62 11.575 3.04 11.805 3.04 11.805 3.62 13.47 3.62 13.765 3.62 13.765 3.04 13.995 3.04 13.995 3.62 14.56 3.62 14.56 4.22 13.47 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 14.095 0.3 14.095 0.83 13.865 0.83 13.865 0.3 11.855 0.3 11.855 0.83 11.625 0.83 11.625 0.3 9.49 0.3 9.49 0.655 9.15 0.655 9.15 0.3 7.195 0.3 7.195 0.71 6.965 0.71 6.965 0.3 4.955 0.3 4.955 0.71 4.725 0.71 4.725 0.3 2.715 0.3 2.715 0.71 2.485 0.71 2.485 0.3 0.53 0.3 0.53 0.655 0.19 0.655 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.67 3.16 8.78 3.16 8.78 1.88 9.195 1.88 9.195 1.17 6.505 1.17 6.505 0.76 5.415 0.76 5.415 1.17 4.26 1.17 4.26 0.76 3.175 0.76 3.175 1.17 1.31 1.17 1.31 0.53 1.65 0.53 1.65 0.94 2.945 0.94 2.945 0.53 4.49 0.53 4.49 0.94 5.185 0.94 5.185 0.53 6.735 0.53 6.735 0.94 8.03 0.94 8.03 0.53 8.37 0.53 8.37 0.94 9.425 0.94 9.425 1.79 13.47 1.79 13.47 2.13 9.04 2.13 9.04 3.39 4.67 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_4
