# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.93 1.2 3.355 1.2 3.355 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.48 2.165 20.065 2.165 20.72 2.165 20.72 1.15 18.425 1.15 18.425 0.73 18.765 0.73 18.765 0.92 20.72 0.92 20.72 0.675 21.19 0.675 21.19 3.38 20.72 3.38 20.72 2.395 20.065 2.395 18.71 2.395 18.71 3.38 18.48 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.285 12.085 3.285 12.085 3.62 13.395 3.62 17.46 3.62 17.46 2.53 17.69 2.53 17.69 3.62 19.525 3.62 19.525 2.625 19.865 2.625 19.865 3.62 20.065 3.62 21.74 3.62 21.74 2.53 21.97 2.53 21.97 3.62 22.4 3.62 22.4 4.22 20.065 4.22 13.395 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.07 0.3 22.07 0.69 21.84 0.69 21.84 0.3 19.83 0.3 19.83 0.69 19.6 0.69 19.6 0.3 17.41 0.3 17.41 0.69 17.18 0.69 17.18 0.3 12.285 0.3 12.285 0.635 11.945 0.635 11.945 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.33 1.465 5.33 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 5.56 2.875 5.56 1 4.485 1 4.485 0.77 5.79 0.77 5.79 1.52 8.115 1.52 8.115 1.75 5.79 1.75 5.79 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.465 10.61 1.465 10.61 1.805 9.13 1.805 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.665 2.875 10.84 2.875 10.84 1 9.765 1 9.765 0.77 11.07 0.77 11.07 1.52 13.395 1.52 13.395 1.75 11.07 1.75 11.07 3.105 9.665 3.105  ;
        POLYGON 14.18 0.715 14.41 0.715 14.41 1.535 16.36 1.535 16.36 1.875 14.41 1.875 14.41 2.82 14.565 2.82 14.565 3.16 14.18 3.16  ;
        POLYGON 15 2.235 16.65 2.235 16.65 1 14.945 1 14.945 0.77 16.88 0.77 16.88 1.59 20.065 1.59 20.065 1.82 16.88 1.82 16.88 2.465 15.23 2.465 15.23 3.16 15 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_4
