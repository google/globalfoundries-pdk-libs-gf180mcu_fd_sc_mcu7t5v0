# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.16 1.17 5.5 1.17 5.5 1.77 6.11 1.77 6.11 2.15 5.16 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.17 4.39 1.17 4.39 2.135 4.01 2.135  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 1.345 2.11 1.345 2.11 1.575 1.56 1.575 1.56 3.32 1.24 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.345 1 1.345 1 3.32 0.705 3.32  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9645 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 1.21 2.715 1.21 2.945 1.21 2.945 0.61 3.26 0.61 3.26 1.665 2.715 1.665 2.34 1.665  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7536 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.91 2.38 6.11 2.38 6.11 2.93 5.77 2.93 5.77 2.7 4.795 2.7 4.795 2.595 2.77 2.595 2.77 2.93 2.43 2.93 2.43 2.365 4.62 2.365 4.62 0.61 5.095 0.61 5.095 0.91 4.91 0.91  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 3.61 3.62 3.61 3.285 3.95 3.285 3.95 3.62 6.57 3.62 6.72 3.62 6.72 4.22 6.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.625 0.475 0.625 0.475 0.865 1.88 0.865 1.88 0.625 2.715 0.625 2.715 0.965 2.11 0.965 2.11 1.095 0.245 1.095  ;
        POLYGON 2.18 3.16 3.13 3.16 3.13 2.825 4.52 2.825 4.52 3.16 6.34 3.16 6.34 0.91 5.87 0.91 5.87 0.68 6.57 0.68 6.57 3.39 4.29 3.39 4.29 3.055 3.36 3.055 3.36 3.39 1.95 3.39 1.95 1.905 3.54 1.905 3.54 0.68 3.95 0.68 3.95 0.91 3.77 0.91 3.77 2.135 2.18 2.135  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_1
