# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.71 1.21 3.83 1.21 3.83 1.34 7.935 1.34 7.935 1.57 1.71 1.57  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.44 1.8 9.035 1.8 9.035 2.12 1.44 2.12  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.55 1.8 10.57 1.8 10.57 2.36 13.53 2.36 13.53 1.965 13.87 1.965 13.87 2.36 15.205 2.36 15.205 1.965 15.545 1.965 15.545 2.36 18.57 2.36 18.57 1.8 19.59 1.8 19.59 2.12 18.8 2.12 18.8 2.595 10.34 2.595 10.34 2.12 9.55 2.12  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.84 1.505 18.25 1.505 18.25 2.13 16.08 2.13 16.08 1.735 10.84 1.735  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.2952 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.98 0.955 1.19 0.955 1.19 0.7 2.9 0.7 2.9 0.53 3.24 0.53 3.24 0.7 4.71 0.7 4.71 0.87 6.98 0.87 6.98 0.575 7.32 0.575 7.32 0.87 8.735 0.87 8.735 1.045 10.36 1.045 10.36 0.775 10.7 0.775 10.7 1.045 13.04 1.045 13.04 0.775 13.38 0.775 13.38 1.045 15.72 1.045 15.72 0.775 16.06 0.775 16.06 1.045 18.4 1.045 18.4 0.775 18.74 0.775 18.74 1.275 8.505 1.275 8.505 1.1 4.48 1.1 4.48 0.93 1.42 0.93 1.42 1.185 1.21 1.185 1.21 2.36 8.34 2.36 8.34 2.68 0.98 2.68  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 11.7 3.62 11.7 3.285 12.04 3.285 12.04 3.62 16.975 3.62 16.975 3.285 17.315 3.285 17.315 3.62 19.755 3.62 20.16 3.62 20.16 4.22 19.755 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.805 0.3 19.805 1.06 19.575 1.06 19.575 0.3 17.4 0.3 17.4 0.765 17.06 0.765 17.06 0.3 14.72 0.3 14.72 0.765 14.38 0.765 14.38 0.3 12.04 0.3 12.04 0.71 11.7 0.71 11.7 0.3 9.36 0.3 9.36 0.765 9.02 0.765 9.02 0.3 5.28 0.3 5.28 0.64 4.94 0.64 4.94 0.3 0.96 0.3 0.96 0.71 0.62 0.71 0.62 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.86 3.16 9.07 3.16 9.07 2.53 9.41 2.53 9.41 2.825 19.525 2.825 19.525 2.53 19.755 2.53 19.755 3.38 19.525 3.38 19.525 3.055 9.41 3.055 9.41 3.39 0.86 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_4
