# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 7 1.565 7 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.53 2.53 11.65 2.53 11.9 2.53 11.9 1.12 11.31 1.12 11.31 0.6 12.22 0.6 12.22 3.38 11.65 3.38 11.53 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 8.115 3.62 10.51 3.62 10.51 2.815 10.85 2.815 10.85 3.62 11.65 3.62 12.605 3.62 12.605 2.53 12.835 2.53 12.835 3.62 13.44 3.62 13.44 4.22 11.65 4.22 8.115 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 12.935 0.3 12.935 1.075 12.705 1.075 12.705 0.3 10.515 0.3 10.515 1.075 10.285 1.075 10.285 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.775 2.825 7.775 2.25 8.115 2.25 8.115 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.17 1.105 8.17 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.315 2.195 7.315 1.79 8.445 1.79 8.445 0.55 8.675 0.55 8.675 1.79 9.89 1.79 9.89 2.02 8.575 2.02 8.575 3.39 8.345 3.39 8.345 2.02 7.545 2.02 7.545 2.535 6.165 2.535  ;
        POLYGON 9.165 2.34 10.345 2.34 10.345 1.545 9.165 1.545 9.165 0.735 9.395 0.735 9.395 1.315 10.575 1.315 10.575 1.69 11.65 1.69 11.65 2.03 10.575 2.03 10.575 2.57 9.395 2.57 9.395 3.25 9.165 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_2
