# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 6.245 3.62 6.245 2.49 6.475 2.49 6.475 3.62 8.485 3.62 8.485 2.49 8.715 2.49 8.715 3.62 10.725 3.62 10.725 2.49 10.955 2.49 10.955 3.62 12.965 3.62 12.965 2.49 13.195 2.49 13.195 3.62 15.205 3.62 15.205 2.49 15.435 2.49 15.435 3.62 17.445 3.62 17.445 2.49 17.675 2.49 17.675 3.62 17.92 3.62 17.92 4.22 17.675 4.22 15.435 4.22 13.195 4.22 10.955 4.22 8.715 4.22 6.475 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.155 0.3 16.155 1.045 15.925 1.045 15.925 0.3 13.915 0.3 13.915 1.045 13.685 1.045 13.685 0.3 11.675 0.3 11.675 1.045 11.445 1.045 11.445 0.3 9.435 0.3 9.435 1.045 9.205 1.045 9.205 0.3 7.195 0.3 7.195 1.045 6.965 1.045 6.965 0.3 4.955 0.3 4.955 1.045 4.725 1.045 4.725 0.3 2.715 0.3 2.715 1.045 2.485 1.045 2.485 0.3 0.475 0.3 0.475 1.045 0.245 1.045 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
        POLYGON 4.725 1.325 6 1.325 6 1.555 4.955 1.555 4.955 3.39 4.725 3.39  ;
        POLYGON 5.21 1.96 6.245 1.96 6.245 0.53 6.475 0.53 6.475 2.19 5.21 2.19  ;
        POLYGON 6.965 1.325 8.24 1.325 8.24 1.555 7.195 1.555 7.195 3.39 6.965 3.39  ;
        POLYGON 7.45 1.96 8.485 1.96 8.485 0.53 8.715 0.53 8.715 2.19 7.45 2.19  ;
        POLYGON 9.205 1.325 10.48 1.325 10.48 1.555 9.435 1.555 9.435 3.39 9.205 3.39  ;
        POLYGON 9.69 1.96 10.725 1.96 10.725 0.53 10.955 0.53 10.955 2.19 9.69 2.19  ;
        POLYGON 11.445 1.325 12.72 1.325 12.72 1.555 11.675 1.555 11.675 3.39 11.445 3.39  ;
        POLYGON 11.93 1.96 12.965 1.96 12.965 0.53 13.195 0.53 13.195 2.19 11.93 2.19  ;
        POLYGON 13.685 1.325 14.96 1.325 14.96 1.555 13.915 1.555 13.915 3.39 13.685 3.39  ;
        POLYGON 14.17 1.96 15.205 1.96 15.205 0.53 15.435 0.53 15.435 2.19 14.17 2.19  ;
        POLYGON 15.925 1.325 17.2 1.325 17.2 1.555 16.155 1.555 16.155 3.39 15.925 3.39  ;
        POLYGON 16.41 1.96 17.445 1.96 17.445 0.53 17.675 0.53 17.675 2.19 16.41 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_32
