# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.369 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.745 4.13 1.745 4.13 2.15 0.65 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.99 2.36 12.975 2.36 12.975 3.39 12.745 3.39 12.745 2.68 10.735 2.68 10.735 3.39 10.505 3.39 10.505 2.68 8.92 2.68 8.495 2.68 8.495 3.39 8.265 3.39 8.265 2.68 6.255 2.68 6.255 3.39 6.025 3.39 6.025 2.36 8.92 2.36 9.61 2.36 9.61 1.51 6.025 1.51 6.025 0.69 6.255 0.69 6.255 1.22 8.265 1.22 8.265 0.69 8.495 0.69 8.495 1.22 10.505 1.22 10.505 0.69 10.735 0.69 10.735 1.22 12.745 1.22 12.745 0.69 12.975 0.69 12.975 1.51 9.99 1.51  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.485 3.62 2.485 3.05 2.715 3.05 2.715 3.62 4.905 3.62 4.905 3.23 5.135 3.23 5.135 3.62 7.145 3.62 7.145 3.05 7.375 3.05 7.375 3.62 8.92 3.62 9.385 3.62 9.385 3.05 9.615 3.05 9.615 3.62 11.625 3.62 11.625 3.05 11.855 3.05 11.855 3.62 13.72 3.62 13.865 3.62 13.865 2.76 14.095 2.76 14.095 3.62 14.56 3.62 14.56 4.22 13.72 4.22 8.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.985 9.33 0.985 9.33 0.3 7.43 0.3 7.43 0.985 7.09 0.985 7.09 0.3 5.19 0.3 5.19 1.055 4.85 1.055 4.85 0.3 2.77 0.3 2.77 1.04 2.43 1.04 2.43 0.3 0.53 0.3 0.53 1.04 0.19 1.04 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 4.425 2.53 4.425 1.5 1.365 1.5 1.365 0.74 1.595 0.74 1.595 1.27 3.605 1.27 3.605 0.74 3.835 0.74 3.835 1.27 4.655 1.27 4.655 1.74 8.92 1.74 8.92 1.975 4.655 1.975 4.655 2.76 3.835 2.76 3.835 3.39 3.605 3.39 3.605 2.76 1.595 2.76 1.595 3.39 1.365 3.39  ;
        POLYGON 10.53 1.74 13.72 1.74 13.72 2.04 10.53 2.04  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
