# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 39.2 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.13 1.77 9.85 1.77 9.85 2.15 5.13 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.205 ;
    PORT
      LAYER METAL1 ;
        POLYGON 29.85 2.425 37.785 2.425 37.785 3.38 37.5 3.38 37.5 3.005 35.455 3.005 35.455 3.38 35.225 3.38 35.225 3.005 33.205 3.005 33.205 3.38 32.975 3.38 32.975 3.005 30.985 3.005 30.985 3.38 30.755 3.38 30.755 3.005 28.74 3.005 28.74 3.38 28.51 3.38 28.51 3.005 28.145 3.005 26.485 3.005 26.485 3.38 26.255 3.38 26.255 3.005 24.255 3.005 24.255 3.38 24.025 3.38 24.025 3.005 22.05 3.005 22.05 3.38 21.82 3.38 21.82 2.425 28.145 2.425 28.95 2.425 28.95 1.445 25.24 1.445 25.24 1.135 21.755 1.135 21.755 0.865 37.785 0.865 37.785 1.135 34.285 1.135 34.285 1.445 29.85 1.445  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.63 3.62 1.63 3.285 1.97 3.285 1.97 3.62 5.045 3.62 5.045 3.445 5.385 3.445 5.385 3.62 8.155 3.62 8.155 3.445 8.515 3.445 8.515 3.62 11.35 3.62 11.35 2.7 11.58 2.7 11.58 3.62 13.76 3.62 13.76 2.7 13.99 2.7 13.99 3.62 15.995 3.62 15.995 2.7 16.225 2.7 16.225 3.62 18.33 3.62 18.33 2.7 18.56 2.7 18.56 3.62 20.68 3.62 20.68 2.7 20.91 2.7 20.91 3.62 22.835 3.62 22.835 3.285 23.175 3.285 23.175 3.62 25.08 3.62 25.08 3.285 25.42 3.285 25.42 3.62 27.33 3.62 27.33 3.285 27.67 3.285 27.67 3.62 28.145 3.62 29.57 3.62 29.57 3.285 29.91 3.285 29.91 3.62 31.81 3.62 31.81 3.285 32.15 3.285 32.15 3.62 34.05 3.62 34.05 3.285 34.39 3.285 34.39 3.62 36.285 3.62 36.285 3.285 36.625 3.285 36.625 3.62 38.3 3.62 38.52 3.62 38.52 2.53 38.75 2.53 38.75 3.62 39.2 3.62 39.2 4.22 38.3 4.22 28.145 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 39.2 -0.3 39.2 0.3 38.85 0.3 38.85 1.015 38.62 1.015 38.62 0.3 36.665 0.3 36.665 0.635 36.325 0.635 36.325 0.3 34.425 0.3 34.425 0.635 34.085 0.635 34.085 0.3 32.185 0.3 32.185 0.635 31.845 0.635 31.845 0.3 29.945 0.3 29.945 0.635 29.605 0.635 29.605 0.3 27.705 0.3 27.705 0.635 27.365 0.635 27.365 0.3 25.465 0.3 25.465 0.635 25.125 0.635 25.125 0.3 23.225 0.3 23.225 0.635 22.885 0.635 22.885 0.3 20.93 0.3 20.93 0.87 20.7 0.87 20.7 0.3 18.51 0.3 18.51 0.87 18.28 0.87 18.28 0.3 16.27 0.3 16.27 0.87 16.04 0.87 16.04 0.3 14.03 0.3 14.03 0.87 13.8 0.87 13.8 0.3 11.635 0.3 11.635 0.475 11.275 0.475 11.275 0.3 8.515 0.3 8.515 0.475 8.155 0.475 8.155 0.3 5.385 0.3 5.385 0.53 5.1 0.53 5.1 0.3 1.7 0.3 1.7 0.76 1.47 0.76 1.47 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.665 2.57 2.045 2.57 2.045 1.225 0.35 1.225 0.35 0.675 0.58 0.675 0.58 0.99 2.275 0.99 2.275 2.035 3.375 2.035 3.375 2.8 0.895 2.8 0.895 3.38 0.665 3.38  ;
        POLYGON 6.31 2.525 10.175 2.525 10.175 1.42 6.595 1.42 6.595 0.99 6.955 0.99 6.955 1.19 9.715 1.19 9.715 0.99 10.415 0.99 10.415 1.63 20.325 1.63 20.325 1.96 10.405 1.96 10.405 2.78 9.315 2.78 9.315 2.755 7.125 2.755 7.125 2.78 6.31 2.78  ;
        POLYGON 2.59 0.53 4.87 0.53 4.87 0.76 6.135 0.76 6.135 0.53 7.415 0.53 7.415 0.73 9.255 0.73 9.255 0.53 11.045 0.53 11.045 0.73 13.255 0.73 13.255 1.1 14.92 1.1 14.92 0.53 15.15 0.53 15.15 1.1 17.16 1.1 17.16 0.53 17.39 0.53 17.39 1.1 19.58 1.1 19.58 0.53 19.81 0.53 19.81 1.1 20.93 1.1 20.93 1.365 24.785 1.365 24.785 1.595 20.7 1.595 20.7 1.33 13.025 1.33 13.025 0.96 10.815 0.96 10.815 0.76 9.485 0.76 9.485 0.96 7.185 0.96 7.185 0.76 6.365 0.76 6.365 0.99 4.64 0.99 4.64 0.76 3.31 0.76 3.31 1.575 3.955 1.575 3.955 2.89 3.725 2.89 3.725 1.805 3.08 1.805 3.08 0.885 2.59 0.885  ;
        POLYGON 2.59 3.12 4.185 3.12 4.185 1.345 3.865 1.345 3.865 0.99 4.225 0.99 4.225 1.115 4.415 1.115 4.415 2.985 5.845 2.985 5.845 3.01 7.385 3.01 7.385 2.985 9.085 2.985 9.085 3.01 10.815 3.01 10.815 2.19 20.7 2.19 20.7 1.96 28.145 1.96 28.145 2.195 20.93 2.195 20.93 2.425 19.75 2.425 19.75 3.38 19.52 3.38 19.52 2.425 17.355 2.425 17.355 3.38 17.125 3.38 17.125 2.425 15.11 2.425 15.11 3.38 14.88 3.38 14.88 2.425 12.86 2.425 12.86 3.38 12.63 3.38 12.63 2.425 11.045 2.425 11.045 3.355 8.855 3.355 8.855 3.215 7.615 3.215 7.615 3.355 5.615 3.355 5.615 3.215 4.815 3.215 4.815 3.35 2.59 3.35  ;
        POLYGON 34.765 1.365 38.3 1.365 38.3 1.595 34.765 1.595  ;
        POLYGON 32.315 1.96 38.3 1.96 38.3 2.195 32.315 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_16
