# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.825 0.55 2.12 0.55 2.12 2.135 1.825 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 0.55 1 0.55 1 2.23 0.705 2.23  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.36 1.16 2.66 1.16 2.66 1.8 3.37 1.8 3.37 2.12 2.36 2.12  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.89 1.24 3.94 1.24 3.94 1.8 4.97 1.8 4.97 2.12 3.65 2.12 3.65 1.56 2.89 1.56  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.67285 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.24 0.55 1.595 0.55 1.595 2.365 4.92 2.365 4.92 2.93 4.58 2.93 4.58 2.595 2.77 2.595 2.77 2.93 2.43 2.93 2.43 2.7 1.24 2.7  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.92 0.525 2.92 0.525 3.62 3.55 3.62 3.55 3.285 3.89 3.285 3.89 3.62 5.45 3.62 5.6 3.62 5.6 4.22 5.45 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 0.89 4.725 0.89 4.725 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.55 0.475 0.55 0.475 2.46 0.985 2.46 0.985 3.16 3.06 3.16 3.06 2.825 4.35 2.825 4.35 3.16 5.22 3.16 5.22 1.37 4.24 1.37 4.24 0.835 2.43 0.835 2.43 0.605 4.24 0.605 4.24 0.6 4.47 0.6 4.47 1.14 5.45 1.14 5.45 3.39 4.12 3.39 4.12 3.055 3.29 3.055 3.29 3.39 0.755 3.39 0.755 2.69 0.245 2.69  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_1
