# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.55 1.41 12.18 1.41 12.18 1.64 9.96 1.64 9.96 2.85 9.55 2.85  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.405 1.75 1.57 1.75 1.57 1.87 7.97 1.87 7.97 1.75 9.03 1.75 9.03 2.15 0.405 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 1.41 3.47 1.41 3.47 1.01 3.91 1.01 3.91 1.41 5.7 1.41 5.7 1.01 6.15 1.01 6.15 1.41 7.735 1.41 7.735 1.64 1.79 1.64  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9636 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.19 1.875 12.42 1.875 12.42 1.18 6.45 1.18 6.45 0.76 5.47 0.76 5.47 1.18 4.21 1.18 4.21 0.76 3.23 0.76 3.23 1.18 1.255 1.18 1.255 0.53 1.65 0.53 1.65 0.945 3 0.945 3 0.53 4.44 0.53 4.44 0.945 5.24 0.945 5.24 0.53 6.68 0.53 6.68 0.945 7.95 0.945 7.95 0.53 8.82 0.53 8.82 0.945 9.72 0.945 9.72 0.53 11.16 0.53 11.16 0.945 12.46 0.945 12.46 0.53 12.85 0.53 12.85 2.91 12.46 2.91 12.46 2.11 10.555 2.11 10.555 2.91 10.19 2.91  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.385 3.62 2.385 3.155 2.615 3.155 2.615 3.62 6.865 3.62 6.865 3.155 7.095 3.155 7.095 3.62 13.815 3.62 14.56 3.62 14.56 4.22 13.815 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.97 0.3 13.97 0.655 13.63 0.655 13.63 0.3 11.73 0.3 11.73 0.655 11.39 0.655 11.39 0.3 9.49 0.3 9.49 0.655 9.15 0.655 9.15 0.3 7.25 0.3 7.25 0.655 6.91 0.655 6.91 0.3 5.01 0.3 5.01 0.655 4.67 0.655 4.67 0.3 2.77 0.3 2.77 0.655 2.43 0.655 2.43 0.3 0.53 0.3 0.53 0.655 0.19 0.655 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 2.57 8.22 2.57 8.22 3.16 11.345 3.16 11.345 2.53 11.575 2.53 11.575 3.16 13.585 3.16 13.585 2.53 13.815 2.53 13.815 3.39 7.99 3.39 7.99 2.8 4.855 2.8 4.855 3.38 4.625 3.38 4.625 2.8 0.475 2.8 0.475 3.38 0.245 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor3_4
