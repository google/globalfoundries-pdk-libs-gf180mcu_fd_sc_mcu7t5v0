# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.265 4.905 1.265 4.905 1.535 1.935 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 2.385 3.57 2.385 3.935 2.385 3.935 1.815 5.715 1.815 5.715 2.1 4.24 2.1 4.24 2.655 3.57 2.655 0.825 2.655  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.3 1.815 9.905 1.815 10.17 1.815 10.17 1.21 11.075 1.21 11.075 1.61 10.425 1.61 10.425 2.095 9.905 2.095 8.3 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.015 2.36 14.915 2.36 15.155 2.36 15.155 1.56 12.965 1.56 12.965 0.6 13.31 0.6 13.31 1.24 15.155 1.24 15.155 0.6 15.535 0.6 15.535 3.39 15.155 3.39 15.155 2.68 14.915 2.68 13.295 2.68 13.295 3.39 13.015 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.42 3.62 2.42 2.895 2.78 2.895 2.78 3.62 3.57 3.62 6.055 3.62 9.09 3.62 9.09 2.785 9.43 2.785 9.43 3.62 12.575 3.62 14.035 3.62 14.035 2.95 14.265 2.95 14.265 3.62 14.915 3.62 15.68 3.62 15.68 4.22 14.915 4.22 12.575 4.22 6.055 4.22 3.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 14.315 0.3 14.315 0.975 14.085 0.975 14.085 0.3 12.49 0.3 12.49 0.635 12.15 0.635 12.15 0.3 9.275 0.3 9.275 0.89 9.045 0.89 9.045 0.3 6.91 0.3 6.91 0.76 6.57 0.76 6.57 0.3 6.11 0.3 6.11 0.76 5.77 0.76 5.77 0.3 2.855 0.3 2.855 0.76 2.515 0.76 2.515 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 1.765 3.57 1.765 3.57 1.995 1.365 1.995 1.365 1.225 0.575 1.225 0.575 3.19 0.345 3.19  ;
        POLYGON 3.72 2.895 4.08 2.895 4.08 3.155 5.76 3.155 5.76 2.84 6.055 2.84 6.055 3.39 3.72 3.39  ;
        POLYGON 6.745 1.86 7.69 1.86 7.69 0.53 8.03 0.53 8.03 1.15 9.905 1.15 9.905 1.555 9.515 1.555 9.515 1.38 8.03 1.38 8.03 2.095 7.085 2.095 7.085 2.925 6.745 2.925  ;
        POLYGON 6.515 3.155 7.835 3.155 7.835 2.325 10.655 2.325 10.655 2.24 11.765 2.24 11.765 1.715 11.995 1.715 11.995 2.47 10.885 2.47 10.885 2.555 8.065 2.555 8.065 3.39 6.285 3.39 6.285 2.565 5.09 2.565 5.09 2.925 4.75 2.925 4.75 2.335 6.285 2.335 6.285 1.22 5.23 1.22 5.23 0.76 3.73 0.76 3.73 0.53 5.46 0.53 5.46 0.99 7.435 0.99 7.435 1.225 6.515 1.225  ;
        POLYGON 10.045 3.16 12.575 3.16 12.575 3.39 10.045 3.39  ;
        POLYGON 11.115 2.7 12.345 2.7 12.345 1.095 11.405 1.095 11.405 0.765 10.035 0.765 10.035 0.53 11.71 0.53 11.71 0.865 12.575 0.865 12.575 1.815 14.915 1.815 14.915 2.045 12.575 2.045 12.575 2.93 11.115 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_2
