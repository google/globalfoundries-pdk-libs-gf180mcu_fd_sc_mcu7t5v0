# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__tieh
  CLASS core TIEHIGH ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__tieh 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.5368 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.22 2.305 1.58 2.305 1.58 3.39 1.22 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.25 3.62 0.25 2.36 0.48 2.36 0.48 3.62 1.6 3.62 2.24 3.62 2.24 4.22 1.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.48 0.3 0.48 1.16 0.25 1.16 0.25 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.875 1.335 1.37 1.335 1.37 0.53 1.6 0.53 1.6 1.57 0.875 1.57  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__tieh
