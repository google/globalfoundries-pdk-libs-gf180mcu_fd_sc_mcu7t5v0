* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24 net_7 net_9 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55 net_6 net_8 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27 net_17 net_14 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63 net_16 net_15 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22 net_13 net_11 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93 net_12 net_10 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33 VDD net_7 net_9 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23 VDD net_6 net_8 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94 VDD net_17 net_14 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87 VDD net_16 net_15 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95 VDD net_13 net_11 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23 VDD net_12 net_10 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS
