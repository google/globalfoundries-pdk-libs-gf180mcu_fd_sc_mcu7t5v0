# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.12 1.77 0.63 1.77 0.63 1.03 1 1.03 1 2.15 0.12 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 1.77 1.75 1.77 1.75 1.03 2.12 1.03 2.12 2.15 1.23 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.77 2.87 1.77 2.87 1.03 3.24 1.03 3.24 2.15 2.35 2.15  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 1.77 4.595 1.77 4.595 2.15 3.47 2.15  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.495 0.805 6.07 0.805 6.07 3.235 5.495 3.235  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.3 3.62 0.3 3.16 0.53 3.16 0.53 3.62 2.285 3.62 2.285 3.28 2.625 3.28 2.625 3.62 4.325 3.62 4.325 3.285 4.665 3.285 4.665 3.62 5.23 3.62 6.6 3.62 6.6 2.65 6.83 2.65 6.83 3.62 7.28 3.62 7.28 4.22 5.23 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 6.85 0.3 6.85 0.765 6.62 0.765 6.62 0.3 4.665 0.3 4.665 0.635 4.325 0.635 4.325 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 2.79 5 2.79 5 1.095 3.845 1.095 3.845 0.78 0.235 0.78 0.235 0.55 4.075 0.55 4.075 0.865 5.23 0.865 5.23 3.02 1.26 3.02  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_2
