# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.95 1.265 4.2 1.265 4.2 1.555 1.95 1.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.785 4.53 1.785 4.53 1.26 6.245 1.26 6.245 1.535 5.05 1.535 5.05 2.02 1.77 2.02  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.78 1.77 1.54 1.77 1.54 2.25 5.69 2.25 5.69 1.785 6.67 1.785 6.67 2.15 6.175 2.15 6.175 2.485 1.265 2.485 1.265 2.15 0.78 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.963 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.43 2.715 5.725 2.715 5.725 2.95 0.13 2.95 0.13 0.865 1.04 0.865 1.04 0.705 3.995 0.705 3.995 0.975 1.37 0.975 1.37 1.1 0.43 1.1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.265 3.62 0.265 3.18 0.495 3.18 0.495 3.62 2.305 3.62 2.305 3.18 2.535 3.18 2.535 3.62 4.345 3.62 4.345 3.18 4.575 3.18 4.575 3.62 6.385 3.62 6.385 2.64 6.615 2.64 6.615 3.62 7.28 3.62 7.28 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 6.615 0.3 6.615 0.9 6.385 0.9 6.385 0.3 0.69 0.3 0.69 0.635 0.35 0.635 0.35 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_2
