# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 23.52 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 22.04 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.765 8.02 1.765 8.02 2.15 0.61 2.15  ;
        POLYGON 14.985 1.765 22.375 1.765 22.375 2.15 14.985 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.38 8.395 2.38 8.395 2.315 11.03 2.315 11.03 1.605 8.415 1.605 8.415 1.535 1.31 1.535 1.31 0.73 1.65 0.73 1.65 0.865 3.605 0.865 3.605 0.675 3.835 0.675 3.835 0.865 5.845 0.865 5.845 0.675 6.075 0.675 6.075 0.865 8.085 0.865 8.085 0.675 8.315 0.675 8.315 0.865 10.325 0.865 10.325 0.675 10.555 0.675 10.555 0.865 12.565 0.865 12.565 0.675 12.795 0.675 12.795 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 0.865 19.285 0.865 19.285 0.675 19.515 0.675 19.515 0.865 21.525 0.865 21.525 0.675 21.755 0.675 21.755 1.535 14.77 1.535 14.77 1.605 11.93 1.605 11.93 2.315 14.665 2.315 14.665 2.38 21.655 2.38 21.655 3.375 21.425 3.375 21.425 3.055 19.415 3.055 19.415 3.375 19.185 3.375 19.185 3.055 17.175 3.055 17.175 3.375 16.945 3.375 16.945 3.055 14.935 3.055 14.935 3.375 14.705 3.375 14.705 3.055 12.695 3.055 12.695 3.375 12.465 3.375 12.465 3.055 10.455 3.055 10.455 3.375 10.225 3.375 10.225 3.055 8.215 3.055 8.215 3.375 7.985 3.375 7.985 3.055 5.975 3.055 5.975 3.375 5.745 3.375 5.745 3.055 3.735 3.055 3.735 3.375 3.505 3.375 3.505 3.055 1.595 3.055 1.595 3.375 1.365 3.375  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.33 3.62 2.33 3.285 2.67 3.285 2.67 3.62 4.57 3.62 4.57 3.285 4.91 3.285 4.91 3.62 6.81 3.62 6.81 3.285 7.15 3.285 7.15 3.62 9.05 3.62 9.05 3.285 9.39 3.285 9.39 3.62 11.29 3.62 11.29 3.285 11.63 3.285 11.63 3.62 13.53 3.62 13.53 3.285 13.87 3.285 13.87 3.62 15.77 3.62 15.77 3.285 16.11 3.285 16.11 3.62 18.01 3.62 18.01 3.285 18.35 3.285 18.35 3.62 20.25 3.62 20.25 3.285 20.59 3.285 20.59 3.62 22.545 3.62 22.545 2.64 22.775 2.64 22.775 3.62 23.52 3.62 23.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 23.52 -0.3 23.52 0.3 22.875 0.3 22.875 1.015 22.645 1.015 22.645 0.3 20.69 0.3 20.69 0.635 20.35 0.635 20.35 0.3 18.45 0.3 18.45 0.635 18.11 0.635 18.11 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.73 0.3 11.73 0.635 11.39 0.635 11.39 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_20
