# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.505 1.77 3.27 1.77 3.27 2.365 5.865 2.365 5.865 1.87 6.095 1.87 6.095 2.595 2.775 2.595 2.775 2.15 1.505 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.725 1.79 5.51 1.79 5.51 2.135 3.725 2.135  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.14 0.65 0.575 0.65 0.575 3.37 0.14 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.975 0.65 9.735 0.65 9.735 3.37 9.405 3.37 9.405 1.68 8.975 1.68  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.23 1.595 3.23 1.595 3.62 3.59 3.62 3.59 3.285 3.93 3.285 3.93 3.62 4.33 3.62 4.33 3.285 4.67 3.285 4.67 3.62 8.205 3.62 8.205 3.075 8.435 3.075 8.435 3.62 9.055 3.62 10.08 3.62 10.08 4.22 9.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 8.49 0.3 8.49 1.035 8.15 1.035 8.15 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 4.23 0.53 7.25 0.53 7.25 1.035 6.91 1.035 6.91 0.76 4.57 0.76 4.57 1.035 4.23 1.035  ;
        POLYGON 1.155 2.77 2.37 2.77 2.37 3.1 3.11 3.1 3.11 2.825 6.415 2.825 6.415 1.74 7.91 1.74 7.91 1.97 6.645 1.97 6.645 3.055 3.34 3.055 3.34 3.33 2.14 3.33 2.14 3 0.925 3 0.925 0.87 3.475 0.87 3.475 0.81 3.85 0.81 3.85 1.1 1.155 1.1  ;
        POLYGON 7.01 3.01 7.12 3.01 7.12 2.375 8.14 2.375 8.14 1.495 5.57 1.495 5.57 0.99 5.91 0.99 5.91 1.265 8.37 1.265 8.37 1.91 9.055 1.91 9.055 2.25 8.37 2.25 8.37 2.61 7.35 2.61 7.35 3.24 7.01 3.24  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_1
