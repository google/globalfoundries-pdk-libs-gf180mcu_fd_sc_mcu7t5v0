* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
M_i_12 I A2 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_13 VSS A1 I VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_16 I3 I2 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_17 VSS A3 I3 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_8 Z I3 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_6 net_2 A3 Z VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_7 VSS I2 net_2 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_14 net_4 A2 I VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_15 VDD A1 net_4 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pmos_5p0 W=5.65e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=5.65e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=5.65e-07 L=5e-07
M_i_18 net_5 I2 I3 VNW pmos_5p0 W=5.65e-07 L=5e-07
M_i_19 VDD A3 net_5 VNW pmos_5p0 W=5.65e-07 L=5e-07
M_i_11 net_3 I3 VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_9 Z A3 net_3 VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_10 net_3 I2 Z VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
