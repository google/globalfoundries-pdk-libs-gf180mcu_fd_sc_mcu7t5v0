# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.825 3.51 1.825 4.225 1.825 4.225 1.23 4.525 1.23 4.525 2.095 3.51 2.095 1.935 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.86 1.81 1.7 1.81 1.7 2.325 3.51 2.325 4.795 2.325 4.795 1.8 6.18 1.8 6.18 2.12 5.025 2.12 5.025 2.68 3.51 2.68 3 2.68 3 2.555 1.425 2.555 1.425 2.1 0.86 2.1  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2436 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.27 2.36 11.275 2.36 11.51 2.36 11.51 1.56 8.27 1.56 8.27 0.655 8.5 0.655 8.5 1.24 10.51 1.24 10.51 0.655 10.74 0.655 10.74 1.24 11.78 1.24 11.78 2.68 11.275 2.68 10.69 2.68 10.69 3.38 10.46 3.38 10.46 2.68 8.5 2.68 8.5 3.38 8.27 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.355 3.62 0.355 2.795 0.695 2.795 0.695 3.62 2.395 3.62 2.395 2.785 2.735 2.785 2.735 3.62 3.51 3.62 6.275 3.62 6.275 2.815 6.615 2.815 6.615 3.62 7.25 3.62 7.25 2.53 7.48 2.53 7.48 3.62 9.34 3.62 9.34 3 9.57 3 9.57 3.62 11.275 3.62 11.53 3.62 11.53 3 11.76 3 11.76 3.62 12.32 3.62 12.32 4.22 11.275 4.22 3.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.86 0.3 11.86 0.985 11.63 0.985 11.63 0.3 9.62 0.3 9.62 0.985 9.39 0.985 9.39 0.3 7.38 0.3 7.38 0.905 7.15 0.905 7.15 0.3 2.915 0.3 2.915 0.76 2.575 0.76 2.575 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.355 0.53 0.695 0.53 0.695 0.99 3.51 0.99 3.51 1.555 3.17 1.555 3.17 1.22 0.585 1.22 0.585 2.33 1.19 2.33 1.19 2.785 1.805 2.785 1.805 3.015 0.93 3.015 0.93 2.565 0.355 2.565  ;
        POLYGON 3.605 0.53 6.725 0.53 6.725 0.76 3.605 0.76  ;
        POLYGON 3.66 2.965 5.45 2.965 5.45 2.35 6.495 2.35 6.495 1.22 4.92 1.22 4.92 0.99 6.725 0.99 6.725 1.815 11.275 1.815 11.275 2.105 6.725 2.105 6.725 2.585 5.68 2.585 5.68 3.195 3.66 3.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_4
