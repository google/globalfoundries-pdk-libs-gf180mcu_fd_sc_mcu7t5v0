# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 30.24 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.1185 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.615 1.77 8.475 1.77 8.475 2.15 4.615 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.594 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.445 2.46 22.65 2.46 23.04 2.46 23.04 1.265 20.75 1.265 20.75 1.135 17.12 1.135 17.12 0.865 28.88 0.865 28.88 1.135 26.61 1.135 26.61 1.265 23.44 1.265 23.44 2.46 28.28 2.46 28.28 3.38 28.045 3.38 28.045 2.86 26.235 2.86 26.235 3.38 26.005 3.38 26.005 2.86 24.195 2.86 24.195 3.38 23.965 3.38 23.965 2.86 22.65 2.86 22.055 2.86 22.055 3.38 21.825 3.38 21.825 2.86 19.815 2.86 19.815 3.38 19.585 3.38 19.585 2.86 17.675 2.86 17.675 3.38 17.445 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.63 3.62 1.63 3.13 1.86 3.13 1.86 3.62 6.4 3.62 6.4 3.445 6.74 3.445 6.74 3.62 9.815 3.62 9.815 3.1 10.045 3.1 10.045 3.62 12.02 3.62 12.02 2.59 12.36 2.59 12.36 3.62 14.06 3.62 14.06 2.59 14.4 2.59 14.4 3.62 16.17 3.62 16.17 2.59 16.51 2.59 16.51 3.62 18.465 3.62 18.465 3.23 18.695 3.23 18.695 3.62 20.705 3.62 20.705 3.23 20.935 3.23 20.935 3.62 22.65 3.62 22.945 3.62 22.945 3.23 23.175 3.23 23.175 3.62 24.985 3.62 24.985 3.23 25.215 3.23 25.215 3.62 27.025 3.62 27.025 3.23 27.255 3.23 27.255 3.62 28.84 3.62 29.065 3.62 29.065 2.53 29.295 2.53 29.295 3.62 29.485 3.62 30.24 3.62 30.24 4.22 29.485 4.22 28.84 4.22 22.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 30.24 -0.3 30.24 0.3 29.945 0.3 29.945 0.915 29.715 0.915 29.715 0.3 27.76 0.3 27.76 0.635 27.225 0.635 27.225 0.3 25.52 0.3 25.52 0.635 25.18 0.635 25.18 0.3 23.28 0.3 23.28 0.635 22.94 0.635 22.94 0.3 21.04 0.3 21.04 0.635 20.7 0.635 20.7 0.3 18.8 0.3 18.8 0.635 18.46 0.635 18.46 0.3 16.505 0.3 16.505 0.93 16.275 0.93 16.275 0.3 14.265 0.3 14.265 0.93 14.035 0.93 14.035 0.3 12.025 0.3 12.025 0.93 11.795 0.93 11.795 0.3 9.63 0.3 9.63 0.475 9.27 0.475 9.27 0.3 6.51 0.3 6.51 0.475 6.15 0.475 6.15 0.3 1.645 0.3 1.645 0.76 1.415 0.76 1.415 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.61 2.57 1.935 2.57 1.935 1.225 0.295 1.225 0.295 0.715 0.525 0.715 0.525 0.99 2.165 0.99 2.165 2.09 3.375 2.09 3.375 2.32 2.165 2.32 2.165 2.865 0.84 2.865 0.84 3.38 0.61 3.38  ;
        POLYGON 5.15 2.525 8.77 2.525 8.77 1.395 4.59 1.395 4.59 0.99 4.95 0.99 4.95 1.165 7.71 1.165 7.71 0.99 8.07 0.99 8.07 1.165 9 1.165 9 1.65 15.965 1.65 15.965 1.9 9 1.9 9 2.78 7.43 2.78 7.43 2.755 5.665 2.755 5.665 2.78 5.15 2.78  ;
        POLYGON 2.535 0.53 5.92 0.53 5.92 0.705 6.925 0.705 6.925 0.53 8.785 0.53 8.785 0.705 11.285 0.705 11.285 1.19 12.915 1.19 12.915 0.58 13.145 0.58 13.145 1.19 15.155 1.19 15.155 0.58 15.385 0.58 15.385 1.19 16.505 1.19 16.505 1.365 20.475 1.365 20.475 1.595 16.275 1.595 16.275 1.42 11.055 1.42 11.055 0.935 8.555 0.935 8.555 0.76 7.155 0.76 7.155 0.935 5.69 0.935 5.69 0.76 3.255 0.76 3.255 1.63 3.9 1.63 3.9 2.89 3.67 2.89 3.67 1.86 3.025 1.86 3.025 0.885 2.535 0.885  ;
        POLYGON 2.595 3.125 4.13 3.125 4.13 1.4 3.81 1.4 3.81 0.99 4.36 0.99 4.36 3.01 5.94 3.01 5.94 2.985 7.2 2.985 7.2 3.01 9.26 3.01 9.26 2.61 11.055 2.61 11.055 2.13 16.275 2.13 16.275 1.96 22.65 1.96 22.65 2.195 16.505 2.195 16.505 2.36 15.365 2.36 15.365 3.38 15.135 3.38 15.135 2.36 13.325 2.36 13.325 3.38 13.095 3.38 13.095 2.36 11.285 2.36 11.285 3.38 11.055 3.38 11.055 2.84 9.49 2.84 9.49 3.355 6.97 3.355 6.97 3.215 6.17 3.215 6.17 3.355 2.595 3.355  ;
        POLYGON 24.405 1.96 28.84 1.96 28.84 2.195 24.405 2.195  ;
        POLYGON 26.86 1.365 29.485 1.365 29.485 1.595 26.86 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_12
