# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.92 1.73 3.83 1.73 3.83 2.15 3.24 2.15 3.24 2.75 2.92 2.75  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.8 1.65 2.12 1.65 2.12 3.31 1.8 3.31  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 1.65 1 1.65 1 3.31 0.705 3.31  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.065 0.61 4.37 0.61 4.37 2.15 4.065 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.185 0.61 5.49 0.61 5.49 2.19 5.185 2.19  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3048 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.47 2.38 4.6 2.38 4.6 0.61 4.955 0.61 4.955 2.7 3.47 2.7  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.59 0.475 2.59 0.475 3.62 5.745 3.62 5.745 3.2 5.975 3.2 5.975 3.62 6.075 3.62 6.72 3.62 6.72 4.22 6.075 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 2.715 0.3 2.715 0.915 2.485 0.915 2.485 0.3 0.475 0.3 0.475 0.915 0.245 0.915 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 2.68 3.05 5.22 3.05 5.22 2.64 5.845 2.64 5.845 0.61 6.075 0.61 6.075 2.87 5.45 2.87 5.45 3.28 2.45 3.28 2.45 1.4 1.365 1.4 1.365 0.61 1.595 0.61 1.595 1.165 3.605 1.165 3.605 0.61 3.835 0.61 3.835 1.4 2.68 1.4  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_1
