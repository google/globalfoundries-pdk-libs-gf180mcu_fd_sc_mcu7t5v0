* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_15 net_9 net_11 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2_26_13 net_16 net_15 net_18 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_3_30_34 net_18 net_15 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2_0_10 net_14 net_16 net_19 VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_3_4_49 net_19 net_16 VSS VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_14 net_6 VPW nmos_5p0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_14 VSS VPW nmos_5p0  W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1_22 net_15 net_9 net_10 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0_35_50 net_17 net_15 VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1_47_46 net_16 net_15 net_17 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0_9_2 net_20 net_16 VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1_22_38 net_14 net_16 net_20 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_14 VDD VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_14 net_5 VNW pmos_5p0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
