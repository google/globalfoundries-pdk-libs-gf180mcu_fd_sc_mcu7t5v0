* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_12 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=8.2e-07 L=6e-07
M_Mn_inv1 VSS I NI VPW nmos_5p0 W=8.2e-07 L=6e-07
M_Mn_inv2 NI I VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_Mn_inv3 VSS I NI VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17_9 VSS NI NI_N VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N NI VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS NI NI_N VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17_10_0 NI_N NI VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn17_9_17_30 VSS NI NI_N VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_89 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1_34 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_49_80 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1_25_35 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_49 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1_25 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_99 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1_33 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_49_88 ZN NI_N VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 VSS NI_N ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pmos_5p0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.095e-06 L=5e-07
M_Mp_inv1 VDD I NI VNW pmos_5p0 W=1.095e-06 L=5e-07
M_Mp_inv2 NI I VDD VNW pmos_5p0 W=1.095e-06 L=5e-07
M_Mp_inv3 VDD I NI VNW pmos_5p0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp14_10 VDD NI NI_P VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp14_11 NI_P NI VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp14_10_8 VDD NI NI_P VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp14_11_21 NI_P NI VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp14_10_8_17 VDD NI NI_P VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_57 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12_96 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_56_105 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12_57_69 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_56 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12_57 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_58 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12_106 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_56_111 ZN NI_P VDD VNW pmos_5p0 W=1.18e-06 L=5e-07
M_mp4_12_57_75 VDD NI_P ZN VNW pmos_5p0 W=1.18e-06 L=5e-07
.ENDS
