# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.64 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.42 1.665 6.745 1.665 6.745 1.45 8.97 1.45 8.97 1.21 9.94 1.21 9.98 1.21 9.98 2.28 9.94 2.28 9.62 2.28 9.62 1.68 6.975 1.68 6.975 1.985 5.42 1.985  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.03 1.77 4.99 1.77 4.99 2.235 7.67 2.235 7.67 1.91 8.35 1.91 8.35 2.69 7.255 2.69 7.255 2.465 4.46 2.465 4.46 2.15 4.03 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.97 1.77 3.8 1.77 3.8 2.695 6.85 2.695 6.85 2.92 9.01 2.92 9.01 1.91 9.24 1.91 9.24 3.26 6.6 3.26 6.6 2.93 3.47 2.93 3.47 2.12 2.97 2.12  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.064 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.28 1.77 2.13 1.77 2.13 2.15 0.28 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.796 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 2.53 2.36 2.53 2.36 0.99 8.6 0.99 8.6 1.22 2.68 1.22 2.68 2.53 3.2 2.53 3.2 3.16 6.35 3.16 6.35 3.39 2.97 3.39 2.97 2.76 1.595 2.76 1.595 3.375 1.365 3.375  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.53 0.525 2.53 0.525 3.62 2.33 3.62 2.33 3.02 2.67 3.02 2.67 3.62 9.49 3.62 9.49 2.53 9.83 2.53 9.83 3.62 9.94 3.62 10.64 3.62 10.64 4.22 9.94 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 10.64 -0.3 10.64 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.18 0.865 1.9 0.865 1.9 0.53 9.94 0.53 9.94 0.76 2.13 0.76 2.13 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_2
