# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 29.68 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.41 1.77 4.43 1.77 4.43 2.15 3.41 2.15  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.816 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0805 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.075 1.21 21.23 1.21 21.23 1.59 20.075 1.59  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6865 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.21 1.77 7.79 1.77 7.79 2.15 6.21 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3055 ;
    PORT
      LAYER METAL1 ;
        POLYGON 25.31 2.055 27.105 2.055 27.44 2.055 27.44 1.345 25.31 1.345 25.31 0.805 25.54 0.805 25.54 1.115 27.44 1.115 27.44 0.595 27.91 0.595 27.91 3.38 27.44 3.38 27.44 2.29 27.105 2.29 25.64 2.29 25.64 3.38 25.31 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.25 3.62 5.25 3.305 5.59 3.305 5.59 3.62 8.1 3.62 8.1 3.35 8.44 3.35 8.44 3.62 10.85 3.62 11.29 3.62 13.51 3.62 13.51 3.36 13.85 3.36 13.85 3.62 15.985 3.62 15.985 2.93 16.215 2.93 16.215 3.62 17.99 3.62 19.93 3.62 19.93 2.66 20.27 2.66 20.27 3.62 21.235 3.62 22.285 3.62 22.285 2.53 22.515 2.53 22.515 3.62 24.325 3.62 24.325 2.53 24.555 2.53 24.555 3.62 26.38 3.62 26.38 2.53 26.61 2.53 26.61 3.62 27.105 3.62 28.57 3.62 28.57 2.53 28.8 2.53 28.8 3.62 29.68 3.62 29.68 4.22 27.105 4.22 21.235 4.22 17.99 4.22 11.29 4.22 10.85 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 29.68 -0.3 29.68 0.3 28.9 0.3 28.9 1.145 28.67 1.145 28.67 0.3 26.715 0.3 26.715 0.75 26.375 0.75 26.375 0.3 24.42 0.3 24.42 1.145 24.19 1.145 24.19 0.3 22.18 0.3 22.18 1.02 21.95 1.02 21.95 0.3 14.19 0.3 14.19 0.915 13.85 0.915 13.85 0.3 8.41 0.3 8.41 0.475 8.07 0.475 8.07 0.3 5.79 0.3 5.79 0.475 5.45 0.475 5.45 0.3 1.595 0.3 1.595 1.16 1.365 1.16 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.6 2.385 2.6 2.105 2.83 2.105 2.83 2.385 4.725 2.385 4.725 1.455 5.065 1.455 5.065 2.615 0.475 2.615 0.475 3.14 0.245 3.14  ;
        POLYGON 6.785 2.43 8.815 2.43 8.815 1.395 6.51 1.395 6.51 0.99 6.85 0.99 6.85 1.165 9.045 1.165 9.045 2.66 7.07 2.66 7.07 2.835 6.785 2.835  ;
        POLYGON 3.27 2.845 6.05 2.845 6.05 3.16 7.56 3.16 7.56 2.89 9.095 2.89 9.095 3.065 10.51 3.065 10.51 2.655 10.85 2.655 10.85 3.295 8.865 3.295 8.865 3.12 7.79 3.12 7.79 3.39 5.82 3.39 5.82 3.075 3.27 3.075  ;
        POLYGON 3.27 0.705 6.02 0.705 6.02 0.53 7.84 0.53 7.84 0.705 9.085 0.705 9.085 0.53 10.895 0.53 10.895 0.97 10.665 0.97 10.665 0.76 9.315 0.76 9.315 0.935 7.61 0.935 7.61 0.76 6.25 0.76 6.25 0.935 3.61 0.935 3.61 1.095 3.27 1.095  ;
        POLYGON 9.395 2.495 9.71 2.495 9.71 0.99 10.05 0.99 10.05 2.045 11.29 2.045 11.29 2.28 9.995 2.28 9.995 2.835 9.395 2.835  ;
        POLYGON 11.585 1.725 11.785 1.725 11.785 0.68 12.015 0.68 12.015 1.725 14.67 1.725 14.67 1.96 11.815 1.96 11.815 3.015 11.585 3.015  ;
        POLYGON 12.31 1.26 14.745 1.26 14.745 0.53 16.81 0.53 16.81 0.76 14.975 0.76 14.975 1.495 12.31 1.495  ;
        POLYGON 12.85 2.19 14.965 2.19 14.965 1.805 16.03 1.805 16.03 0.99 16.37 0.99 16.37 1.805 17.51 1.805 17.51 2.81 17.17 2.81 17.17 2.04 15.25 2.04 15.25 2.78 14.91 2.78 14.91 2.425 12.85 2.425  ;
        POLYGON 12.11 2.9 14.55 2.9 14.55 3.16 15.48 3.16 15.48 2.465 16.93 2.465 16.93 3.04 17.99 3.04 17.99 3.31 16.7 3.31 16.7 2.7 15.71 2.7 15.71 3.39 14.32 3.39 14.32 3.13 12.45 3.13 12.45 3.355 12.11 3.355  ;
        POLYGON 19.495 2.2 21.235 2.2 21.235 2.835 21.005 2.835 21.005 2.43 19.495 2.43 19.495 2.89 19.265 2.89 19.265 1.22 18.27 1.22 18.27 0.99 19.77 0.99 19.77 1.22 19.495 1.22  ;
        POLYGON 17.15 0.99 17.81 0.99 17.81 0.53 21.72 0.53 21.72 1.45 22.775 1.45 22.775 1.685 21.49 1.685 21.49 0.76 18.04 0.76 18.04 1.875 18.475 1.875 18.475 2.89 18.245 2.89 18.245 2.105 17.81 2.105 17.81 1.22 17.15 1.22  ;
        POLYGON 21.53 1.965 23.07 1.965 23.07 0.805 23.3 0.805 23.3 1.575 27.105 1.575 27.105 1.805 23.535 1.805 23.535 3.38 23.305 3.38 23.305 2.195 21.53 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
