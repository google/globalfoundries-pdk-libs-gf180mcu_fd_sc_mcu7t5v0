# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 6.78 1.565 6.78 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.84 1.085 9.4 1.085 9.4 2.355 8.84 2.355  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.38 2.15 12.745 2.15 12.98 2.15 12.98 1.365 12.38 1.365 12.38 0.545 12.76 0.545 12.76 1.135 13.34 1.135 13.34 2.38 12.76 2.38 12.76 3.38 12.745 3.38 12.38 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 7.875 3.62 9.345 3.62 9.345 2.655 9.575 2.655 9.575 3.62 11.21 3.62 11.21 2.63 11.55 2.63 11.55 3.62 12.745 3.62 13.35 3.62 13.35 2.63 13.69 2.63 13.69 3.62 14 3.62 14 4.22 12.745 4.22 7.875 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14 -0.3 14 0.3 13.735 0.3 13.735 0.885 13.505 0.885 13.505 0.3 11.495 0.3 11.495 0.885 11.265 0.885 11.265 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.535 2.825 7.535 2.25 7.875 2.25 7.875 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.095 1.105 8.095 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.03 2.195 7.03 1.79 8.325 1.79 8.325 0.605 9.895 0.605 9.895 1.67 10.985 1.67 10.985 1.9 9.665 1.9 9.665 0.835 8.555 0.835 8.555 3.39 8.325 3.39 8.325 2.02 7.28 2.02 7.28 2.535 6.165 2.535  ;
        POLYGON 10.245 2.15 11.325 2.15 11.325 1.365 10.145 1.365 10.145 0.545 10.375 0.545 10.375 1.135 11.555 1.135 11.555 1.67 12.745 1.67 12.745 1.9 11.555 1.9 11.555 2.38 10.475 2.38 10.475 3.38 10.245 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
