# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.66 1.065 1.02 1.065 1.02 2.24 0.66 2.24  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.515 2.13 1.515 2.13 3.37 1.77 3.37  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0719 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.42 0.55 3.83 0.55 3.83 3.355 3.42 3.355  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.26 3.62 0.26 2.545 0.49 2.545 0.49 3.62 2.52 3.62 2.52 2.53 2.75 2.53 2.75 3.62 3.19 3.62 4.56 3.62 4.56 2.53 4.79 2.53 4.79 3.62 5.04 3.62 5.04 4.22 3.19 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.79 0.3 4.79 0.765 4.56 0.765 4.56 0.3 2.53 0.3 2.53 0.69 2.3 0.69 2.3 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.195 0.55 1.51 0.55 1.51 0.93 3.19 0.93 3.19 1.755 2.96 1.755 2.96 1.165 1.51 1.165 1.51 3.355 1.28 3.355 1.28 0.78 0.195 0.78  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_2
