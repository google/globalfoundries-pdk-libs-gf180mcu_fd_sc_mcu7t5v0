# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.875 1.82 3.51 1.82 3.785 1.82 3.785 1.34 4.525 1.34 4.525 1.57 4.015 1.57 4.015 2.1 3.51 2.1 1.875 2.1  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.88 1.69 1.56 1.69 1.56 2.33 3.51 2.33 4.255 2.33 4.255 1.8 5.49 1.8 5.49 2.155 4.495 2.155 4.495 2.56 3.51 2.56 2.325 2.56 2.325 2.73 0.88 2.73  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.75 2.695 5.72 2.695 5.72 1.11 3.785 1.11 3.785 0.53 4.015 0.53 4.015 0.875 6.04 0.875 6.04 2.925 4.75 2.925  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.71 3.62 2.71 2.79 3.05 2.79 3.05 3.62 3.51 3.62 6.12 3.62 6.72 3.62 6.72 4.22 6.12 4.22 3.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 6.11 0.3 6.11 0.635 5.77 0.635 5.77 0.3 2.95 0.3 2.95 0.76 2.61 0.76 2.61 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.29 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 0.99 3.51 0.99 3.51 1.555 3.17 1.555 3.17 1.29 0.63 1.29 0.63 3.35 0.29 3.35  ;
        POLYGON 3.59 3.155 6.12 3.155 6.12 3.39 3.59 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_1
