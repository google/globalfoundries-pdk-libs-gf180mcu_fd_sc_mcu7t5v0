# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.455 2.225 1.455 2.225 1.825 3.495 1.825 3.67 1.825 3.67 1.455 4.77 1.455 4.77 1.69 3.9 1.69 3.9 2.095 3.495 2.095 1.77 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.385 3.495 2.385 4.13 2.385 4.13 1.92 5.175 1.92 5.175 1.595 5.62 1.595 5.62 2.15 4.36 2.15 4.36 2.655 3.495 2.655 0.87 2.655  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.085 1.825 9.54 1.825 10.765 1.825 10.765 2.095 9.54 2.095 8.085 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5111 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.57 2.92 11.88 2.92 11.88 2.36 12.17 2.36 12.44 2.36 12.44 1.58 11.17 1.58 11.17 0.99 12.76 0.99 12.76 2.68 12.215 2.68 12.215 3.24 12.17 3.24 9.57 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.37 3.62 2.37 2.9 2.73 2.9 2.73 3.62 3.495 3.62 6.12 3.62 6.545 3.62 6.545 2.84 6.775 2.84 6.775 3.62 8.76 3.62 8.76 2.815 9.1 2.815 9.1 3.62 12.17 3.62 12.465 3.62 12.465 3.015 12.695 3.015 12.695 3.62 12.86 3.62 13.44 3.62 13.44 4.22 12.86 4.22 12.17 4.22 6.12 4.22 3.495 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 8.87 0.3 8.87 0.76 8.53 0.76 8.53 0.3 6.11 0.3 6.11 0.76 5.77 0.76 5.77 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 0.99 1.305 0.99 1.305 0.53 1.65 0.53 1.65 0.99 3.495 0.99 3.495 1.22 0.575 1.22 0.575 3.195 0.345 3.195  ;
        POLYGON 3.72 2.9 4.08 2.9 4.08 3.16 5.76 3.16 5.76 2.9 6.12 2.9 6.12 3.39 3.72 3.39  ;
        POLYGON 6.49 0.53 6.83 0.53 6.83 0.99 9.54 0.99 9.54 1.565 9.2 1.565 9.2 1.225 7.85 1.225 7.85 2.93 7.51 2.93 7.51 1.225 6.49 1.225  ;
        POLYGON 4.74 2.38 5.88 2.38 5.88 1.225 3.73 1.225 3.73 0.53 4.07 0.53 4.07 0.99 6.11 0.99 6.11 2.38 7.03 2.38 7.03 1.535 7.26 1.535 7.26 3.16 8.27 3.16 8.27 2.33 11.22 2.33 11.22 1.86 12.17 1.86 12.17 2.095 11.45 2.095 11.45 2.565 8.5 2.565 8.5 3.39 7.03 3.39 7.03 2.61 5.1 2.61 5.1 2.93 4.74 2.93  ;
        POLYGON 9.74 0.53 12.86 0.53 12.86 0.76 9.74 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_1
