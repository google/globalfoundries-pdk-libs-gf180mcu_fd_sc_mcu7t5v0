# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.725 1.78 18.75 1.78 20.415 1.78 20.415 2.12 18.75 2.12 18.725 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.075 1.78 15.975 1.78 15.975 2.13 14.075 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 1.025 1.01 1.025 1.01 2.835 0.705 2.835  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.505 0.55 4.935 0.55 4.935 1.8 5.755 1.8 5.755 2.15 4.505 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.255 1.8 3.3 1.8 3.3 1.24 3.7 1.24 3.7 2.25 2.255 2.25  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.41 1.305 11.775 1.305 11.775 1.77 12.19 1.77 12.775 1.77 12.775 3.32 12.405 3.32 12.405 2.15 12.19 2.15 11.41 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2064 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.23 0.6 6.6 0.6 6.6 1.8 8.425 1.8 8.425 0.6 8.84 0.6 8.84 2.925 8.425 2.925 8.425 2.15 6.615 2.15 6.615 2.925 6.23 2.925  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.575 0.475 2.575 0.475 3.62 1.65 3.62 5.12 3.62 5.12 2.845 5.46 2.845 5.46 3.62 7.35 3.62 7.35 2.845 7.69 2.845 7.69 3.62 9.53 3.62 9.53 2.845 9.87 2.845 9.87 3.62 10.72 3.62 12.19 3.62 15.145 3.62 15.145 2.845 15.49 2.845 15.49 3.62 17.575 3.62 19.43 3.62 19.43 2.815 19.77 2.815 19.77 3.62 20.935 3.62 21.28 3.62 21.28 4.22 20.935 4.22 17.575 4.22 12.19 4.22 10.72 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 19.815 0.3 19.815 1.145 19.585 1.145 19.585 0.3 15.335 0.3 15.335 1.145 15.105 1.145 15.105 0.3 9.875 0.3 9.875 1.16 9.645 1.16 9.645 0.3 7.635 0.3 7.635 1.16 7.405 1.16 7.405 0.3 5.395 0.3 5.395 1.16 5.165 1.16 5.165 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 2.95 1.26 2.95  ;
        POLYGON 3.93 0.78 4.275 0.78 4.275 2.87 3.93 2.87  ;
        POLYGON 10.335 2.38 10.72 2.38 10.72 3.005 10.49 3.005 10.49 2.615 9.3 2.615 9.3 3.39 7.92 3.39 7.92 2.615 7.12 2.615 7.12 3.39 5.755 3.39 5.755 2.615 4.735 2.615 4.735 3.33 2.71 3.33 2.71 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.91 0.845 2.91 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 3.05 2.74 3.05 3.1 4.505 3.1 4.505 2.38 5.985 2.38 5.985 3.16 6.89 3.16 6.89 2.38 8.15 2.38 8.15 3.155 9.07 3.155 9.07 2.38 10.105 2.38 10.105 0.79 10.72 0.79 10.72 1.13 10.335 1.13  ;
        POLYGON 10.565 1.46 10.95 1.46 10.95 0.845 12.19 0.845 12.19 1.075 11.18 1.075 11.18 2.72 12.12 2.72 12.12 2.95 10.95 2.95 10.95 1.82 10.565 1.82  ;
        POLYGON 13.835 2.575 14.315 2.575 14.315 2.925 13.585 2.925 13.585 0.795 14.315 0.795 14.315 1.145 13.835 1.145  ;
        POLYGON 16.225 0.78 16.455 0.78 16.455 2.925 16.225 2.925  ;
        POLYGON 13.125 0.78 13.355 0.78 13.355 3.16 14.6 3.16 14.6 2.38 15.97 2.38 15.97 3.16 17.245 3.16 17.245 0.78 17.575 0.78 17.575 3.39 15.74 3.39 15.74 2.615 14.83 2.615 14.83 3.39 13.125 3.39  ;
        POLYGON 17.805 0.85 18.75 0.85 18.75 1.08 18.035 1.08 18.035 2.815 18.665 2.815 18.665 3.045 17.805 3.045  ;
        POLYGON 18.265 1.675 18.495 1.675 18.495 2.355 20.705 2.355 20.705 0.78 20.935 0.78 20.935 3.14 20.6 3.14 20.6 2.585 18.265 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_4
