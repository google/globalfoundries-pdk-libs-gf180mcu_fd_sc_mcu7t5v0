* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nmos_5p0 W=3.6e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=4.85e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=4.85e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pmos_5p0 W=1.02e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
