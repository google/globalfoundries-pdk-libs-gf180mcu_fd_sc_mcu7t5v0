# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 1.625 1.59 1.625 1.59 2.125 0.41 2.125  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.082 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.405 1.16 7.77 1.16 7.77 1.64 8.775 1.64 8.775 2.19 7.405 2.19  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.04 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.795 0.53 7.175 0.53 7.175 2.8 6.88 2.8 6.88 1.66 6.795 1.66  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.465 3.62 1.465 2.815 1.805 2.815 1.805 3.62 5.925 3.62 5.925 2.89 6.155 2.89 6.155 3.62 7.965 3.62 7.965 2.98 8.195 2.98 8.195 3.62 9.285 3.62 9.52 3.62 9.52 4.22 9.285 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 8.145 0.3 8.145 0.92 7.915 0.92 7.915 0.3 5.96 0.3 5.96 0.635 5.62 0.635 5.62 0.3 1.605 0.3 1.605 0.76 1.375 0.76 1.375 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.5 2.355 1.84 2.355 1.84 1.225 0.255 1.225 0.255 0.57 0.485 0.57 0.485 0.99 2.07 0.99 2.07 2.035 3.21 2.035 3.21 2.585 0.73 2.585 0.73 3.38 0.5 3.38  ;
        POLYGON 2.495 0.53 5.39 0.53 5.39 0.865 6.565 0.865 6.565 1.64 6.335 1.64 6.335 1.095 5.16 1.095 5.16 0.76 3.215 0.76 3.215 1.575 3.79 1.575 3.79 2.89 3.555 2.89 3.555 1.805 2.985 1.805 2.985 0.885 2.495 0.885  ;
        POLYGON 2.445 3.125 4.02 3.125 4.02 1.345 3.77 1.345 3.77 0.99 4.25 0.99 4.25 1.325 6.105 1.325 6.105 1.965 6.65 1.965 6.65 2.195 5.875 2.195 5.875 1.555 4.25 1.555 4.25 3.125 4.905 3.125 4.905 2.465 5.135 2.465 5.135 3.355 2.445 3.355  ;
        POLYGON 5.415 1.915 5.645 1.915 5.645 2.425 6.615 2.425 6.615 3.07 7.505 3.07 7.505 2.52 9.02 2.52 9.02 0.58 9.285 0.58 9.285 3.38 9.02 3.38 9.02 2.75 7.735 2.75 7.735 3.3 6.385 3.3 6.385 2.66 5.415 2.66  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_2
