# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.76 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.965 1.79 3.27 1.79 3.27 2.12 0.965 2.12  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.78 1.24 4.045 1.24 4.045 2.795 3.5 2.795 3.5 1.56 0.78 1.56  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.38 1.8 7.38 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.895 2.53 11.32 2.53 11.32 1.065 10.75 1.065 10.75 0.6 11.63 0.6 11.63 3.38 10.895 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 2.815 1.55 2.815 1.55 3.62 3.16 3.62 5.365 3.62 5.365 3 5.595 3 5.595 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 10.005 3.62 10.005 2.53 10.235 2.53 10.235 3.62 10.75 3.62 11.76 3.62 11.76 4.22 10.75 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 11.76 -0.3 11.76 0.3 9.955 0.3 9.955 1.075 9.725 1.075 9.725 0.3 5.695 0.3 5.695 0.86 5.465 0.86 5.465 0.3 1.595 0.3 1.595 0.86 1.365 0.86 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 2.35 3.16 2.35 3.16 2.58 0.53 2.58 0.53 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 0.76 3.41 0.76 3.41 0.53 4.56 0.53 4.56 1.225 6.53 1.225 6.53 1.455 4.56 1.455 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.805 9.285 1.805 9.285 2.145 7.97 2.145 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 8.605 2.395 9.525 2.395 9.525 1.555 8.605 1.555 8.605 0.735 8.835 0.735 8.835 1.325 9.755 1.325 9.755 1.79 10.75 1.79 10.75 2.02 9.755 2.02 9.755 2.625 8.835 2.625 8.835 3.25 8.605 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_1
