* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
M_tn9 ncki CLKN VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn16 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 VSS D net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net2 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 ncki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 ncki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn6_7 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp9 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp16 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp10 VDD D net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp11 net5 ncki net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp0 net4 cki net5 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp7 net0 cki net10 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp6 net7 ncki net0 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp2 VDD net1 net7 VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp4_13 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
.ENDS
