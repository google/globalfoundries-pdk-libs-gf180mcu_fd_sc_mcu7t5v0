# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 1.8 13.88 1.8 13.88 2.12 9.57 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 1.76 1.295 1.76 1.295 2.35 4.365 2.35 4.365 1.825 5.725 1.825 5.725 2.35 8.895 2.35 8.895 1.76 9.135 1.76 9.135 2.58 6.365 2.58 6.365 2.69 3.73 2.69 3.73 2.58 1.055 2.58  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 1.8 3.64 1.8 3.64 1.345 6.44 1.345 6.44 1.8 8.35 1.8 8.35 2.12 6.21 2.12 6.21 1.575 3.87 1.575 3.87 2.12 1.73 2.12  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.005 1.8 17.64 1.8 17.64 1.45 20.44 1.45 20.44 1.8 22.35 1.8 22.35 2.12 20.21 2.12 20.21 1.68 17.87 1.68 17.87 2.12 16.005 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 1.8 15.775 1.8 15.775 2.36 18.325 2.36 18.325 1.91 19.685 1.91 19.685 2.36 22.965 2.36 22.965 1.76 23.225 1.76 23.225 2.68 19.945 2.68 19.945 2.595 18.05 2.595 18.05 2.68 15.545 2.68 15.545 2.12 14.65 2.12  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.1761 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 2.36 14.12 2.36 14.12 0.99 22.535 0.99 22.535 1.22 14.42 1.22 14.42 2.36 15.295 2.36 15.295 2.92 18.335 2.92 18.335 2.825 19.655 2.825 19.655 2.92 21.81 2.92 21.81 3.24 19.425 3.24 19.425 3.055 18.585 3.055 18.585 3.24 15.045 3.24 15.045 2.815 9.57 2.815  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.635 3.62 2.635 3.285 2.975 3.285 2.975 3.62 7.115 3.62 7.115 3.285 7.455 3.285 7.455 3.62 14.085 3.62 14.455 3.62 14.455 3.285 14.795 3.285 14.795 3.62 18.835 3.62 18.835 3.285 19.175 3.285 19.175 3.62 23.5 3.62 23.5 2.53 23.73 2.53 23.73 3.62 23.885 3.62 24.08 3.62 24.08 4.22 23.885 4.22 14.085 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 13.055 0.3 13.055 0.635 12.715 0.635 12.715 0.3 10.815 0.3 10.815 0.635 10.475 0.635 10.475 0.3 8.575 0.3 8.575 0.635 8.235 0.635 8.235 0.3 6.335 0.3 6.335 0.635 5.995 0.635 5.995 0.3 4.095 0.3 4.095 0.635 3.755 0.635 3.755 0.3 1.855 0.3 1.855 0.635 1.515 0.635 1.515 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.5 2.53 0.73 2.53 0.73 2.825 3.48 2.825 3.48 2.94 6.615 2.94 6.615 2.825 8.42 2.825 8.42 3.14 14.085 3.14 14.085 3.37 8.19 3.37 8.19 3.055 6.865 3.055 6.865 3.17 3.23 3.17 3.23 3.055 0.73 3.055 0.73 3.38 0.5 3.38  ;
        POLYGON 0.385 0.865 13.405 0.865 13.405 0.53 23.885 0.53 23.885 0.76 13.635 0.76 13.635 1.095 0.385 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_4
