* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_4 Z_neg A1 VDD VNW pfet_05v0 W=6e-07 L=5e-07
M_i_5 VDD A2 Z_neg VNW pfet_05v0 W=6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS
