# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.88 1.24 4.42 1.24 4.42 1.535 1.88 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 1.565 1.105 1.565 1.105 2.265 3.22 2.265 3.45 2.265 3.45 1.82 5.26 1.82 5.26 2.095 3.89 2.095 3.89 2.495 3.22 2.495 0.875 2.495  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5105 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.175 1.8 9.745 1.8 10.02 1.8 10.02 1.255 11.15 1.255 11.15 1.565 10.275 1.565 10.275 2.095 9.745 2.095 8.175 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.94 2.36 17.06 2.36 17.32 2.36 17.32 1.535 12.84 1.535 12.84 0.655 13.07 0.655 13.07 1.26 15.08 1.26 15.08 0.655 15.31 0.655 15.31 1.26 17.32 1.26 17.32 0.6 17.775 0.6 17.775 3.38 17.22 3.38 17.22 2.68 17.06 2.68 15.26 2.68 15.26 3.38 15.03 3.38 15.03 2.68 13.17 2.68 13.17 3.38 12.94 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.33 3.62 2.33 2.725 2.67 2.725 2.67 3.62 3.22 3.62 6.165 3.62 8.965 3.62 8.965 2.785 9.305 2.785 9.305 3.62 12.375 3.62 13.96 3.62 13.96 3.015 14.19 3.015 14.19 3.62 16.15 3.62 16.15 3.015 16.38 3.015 16.38 3.62 17.06 3.62 17.92 3.62 17.92 4.22 17.06 4.22 12.375 4.22 6.165 4.22 3.22 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.43 0.3 16.43 0.905 16.2 0.905 16.2 0.3 14.19 0.3 14.19 0.905 13.96 0.905 13.96 0.3 12.365 0.3 12.365 0.64 12.025 0.64 12.025 0.3 9.145 0.3 9.145 0.84 8.915 0.84 8.915 0.3 6.74 0.3 6.74 0.76 5.59 0.76 5.59 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 1.765 3.22 1.765 3.22 2.035 1.42 2.035 1.42 1.225 0.575 1.225 0.575 3.015 0.345 3.015  ;
        POLYGON 3.55 2.725 3.89 2.725 3.89 3.16 5.825 3.16 5.825 2.725 6.165 2.725 6.165 3.39 3.55 3.39  ;
        POLYGON 6.905 1.8 7.52 1.8 7.52 0.53 7.86 0.53 7.86 1.075 9.745 1.075 9.745 1.56 9.405 1.56 9.405 1.305 7.86 1.305 7.86 2.095 7.245 2.095 7.245 2.93 6.905 2.93  ;
        POLYGON 6.625 3.16 8.115 3.16 8.115 2.325 10.505 2.325 10.505 1.82 11.76 1.82 11.76 2.18 10.735 2.18 10.735 2.555 8.39 2.555 8.39 3.39 6.395 3.39 6.395 2.495 5.67 2.495 5.67 2.555 4.91 2.555 4.91 2.93 4.57 2.93 4.57 2.325 5.44 2.325 5.44 2.265 6.395 2.265 6.395 1.535 5.115 1.535 5.115 0.76 3.55 0.76 3.55 0.53 5.345 0.53 5.345 1.3 7.275 1.3 7.275 1.535 6.625 1.535  ;
        POLYGON 9.895 3.16 12.375 3.16 12.375 3.39 9.895 3.39  ;
        POLYGON 10.915 2.7 12.145 2.7 12.145 1.485 11.565 1.485 11.565 0.76 9.895 0.76 9.895 0.53 11.795 0.53 11.795 1.255 12.375 1.255 12.375 1.765 17.06 1.765 17.06 1.995 12.375 1.995 12.375 2.93 10.915 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_4
