# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.815 1.45 2.22 1.45 2.22 1.825 3.445 1.825 4.57 1.825 4.57 2.095 3.445 2.095 1.815 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.91 1.625 1.535 1.625 1.535 2.385 3.445 2.385 5.185 2.385 5.185 1.51 6.01 1.51 6.01 1.74 5.455 1.74 5.455 2.655 3.445 2.655 1.305 2.655 1.305 1.855 0.91 1.855  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.45635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.305 2.945 3.445 2.945 5.745 2.945 5.745 1.98 6.29 1.98 6.29 1.22 4.98 1.22 4.98 0.99 6.58 0.99 6.58 2.215 6.02 2.215 6.02 3.215 3.445 3.215 3.305 3.215  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.385 3.62 0.385 2.72 0.615 2.72 0.615 3.62 2.65 3.62 2.65 2.93 2.99 2.93 2.99 3.62 3.445 3.62 6.305 3.62 6.305 2.69 6.535 2.69 6.535 3.62 6.69 3.62 7.28 3.62 7.28 4.22 6.69 4.22 3.445 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 2.71 0.3 2.71 0.76 2.37 0.76 2.37 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.33 0.53 0.67 0.53 0.67 0.99 3.445 0.99 3.445 1.565 3.105 1.565 3.105 1.22 0.615 1.22 0.615 2.18 1.075 2.18 1.075 2.945 1.78 2.945 1.78 3.215 0.845 3.215 0.845 2.415 0.33 2.415  ;
        POLYGON 3.63 0.53 6.69 0.53 6.69 0.76 3.63 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_1
