# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.525 1.645 11.06 1.645 11.06 2.365 14.005 2.365 14.005 1.16 14.46 1.16 14.46 2.69 13.285 2.69 13.285 2.595 10.525 2.595  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.29 1.8 13.39 1.8 13.39 2.12 11.29 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.07 2.365 6.04 2.365 6.04 1.79 6.3 1.79 6.3 2.365 9.09 2.365 9.1 2.365 9.1 1.77 9.68 1.77 9.68 2.15 9.38 2.15 9.38 2.595 9.09 2.595 6.74 2.595 6.74 2.69 5.07 2.69  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.77 1.8 8.87 1.8 8.87 2.12 6.77 2.12  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.335 4.38 1.335 4.38 1.8 5.015 1.8 5.015 2.12 4.01 2.12 4.01 1.57 1.02 1.57 1.02 2.19 0.66 2.19  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.8 3.46 1.8 3.46 2.12 1.53 2.12  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.265 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.16 2.825 12.95 2.825 12.95 2.92 14.82 2.92 14.82 3.24 12.72 3.24 12.72 3.055 11.775 3.055 11.775 3.24 9.09 3.24 8.445 3.24 8.445 3.055 7.34 3.055 7.34 3.24 3.125 3.24 3.125 3.055 0.28 3.055 0.28 2.825 3.42 2.825 3.42 2.92 7.09 2.92 7.09 2.825 9.09 2.825 9.93 2.825 9.93 0.99 13.57 0.99 13.57 1.22 10.16 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.285 2.77 3.285 2.77 3.62 7.63 3.62 7.63 3.285 7.97 3.285 7.97 3.62 9.09 3.62 12.11 3.62 12.11 3.285 12.45 3.285 12.45 3.62 14.92 3.62 15.12 3.62 15.12 4.22 14.92 4.22 9.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 0.845 0.245 0.845 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 0.865 5.13 0.865 5.13 0.99 9.09 0.99 9.09 1.22 4.88 1.22 4.88 1.095 1.31 1.095  ;
        POLYGON 5.39 0.53 14.92 0.53 14.92 0.76 5.39 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_2
