# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.605 1.76 4.13 1.76 4.13 2.16 2.605 2.16  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.58 1.76 17.335 1.76 17.335 2.16 16.7 2.16 16.7 3.37 16.34 3.37 16.34 2.16 15.58 2.16  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.754 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.49 1.605 9.695 1.605 14.215 1.605 14.525 1.605 14.525 1.345 14.755 1.345 14.755 1.835 14.215 1.835 9.695 1.835 5.66 1.835 5.66 2.16 4.49 2.16  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0452 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.37 0.55 18.96 0.55 18.96 3.37 18.37 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0062 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.22 0.55 1.68 0.55 1.68 3.37 1.22 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.385 3.62 0.385 2.46 0.615 2.46 0.615 3.62 2.37 3.62 2.37 3.285 2.71 3.285 2.71 3.62 5.83 3.62 7.95 3.62 7.95 3.005 8.29 3.005 8.29 3.62 9.79 3.62 10.53 3.62 10.53 2.845 10.87 2.845 10.87 3.62 12.49 3.62 12.49 3.005 12.83 3.005 12.83 3.62 14.31 3.62 17.405 3.62 17.405 2.48 17.635 2.48 17.635 3.62 18.12 3.62 19.445 3.62 19.445 2.48 19.675 2.48 19.675 3.62 20.16 3.62 20.16 4.22 18.12 4.22 14.31 4.22 9.79 4.22 5.83 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.775 0.3 19.775 0.905 19.545 0.905 19.545 0.3 17.57 0.3 17.57 0.73 17.23 0.73 17.23 0.3 12.93 0.3 12.93 0.915 12.59 0.915 12.59 0.3 10.87 0.3 10.87 1.075 10.53 1.075 10.53 0.3 8.29 0.3 8.29 0.915 7.95 0.915 7.95 0.3 2.755 0.3 2.755 0.695 2.525 0.695 2.525 0.3 0.515 0.3 0.515 0.905 0.285 0.905 0.285 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 2.17 2.61 5.83 2.61 5.83 2.845 1.94 2.845 1.94 0.925 5.545 0.925 5.545 0.78 5.775 0.78 5.775 1.155 2.17 1.155  ;
        POLYGON 6.665 0.79 6.895 0.79 6.895 1.145 9.465 1.145 9.465 0.79 9.695 0.79 9.695 1.375 6.665 1.375  ;
        POLYGON 6.71 2.54 9.79 2.54 9.79 2.775 6.71 2.775  ;
        POLYGON 11.305 0.79 11.535 0.79 11.535 1.145 13.985 1.145 13.985 0.79 14.215 0.79 14.215 1.375 11.305 1.375  ;
        POLYGON 11.24 2.545 14.31 2.545 14.31 2.775 11.24 2.775  ;
        POLYGON 6.07 2.065 15.105 2.065 15.105 0.78 15.335 0.78 15.335 1.085 18.12 1.085 18.12 2.23 17.89 2.23 17.89 1.315 15.335 1.315 15.335 3.14 15.105 3.14 15.105 2.295 6.07 2.295  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_2
