# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.632 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.765 8.51 1.765 8.51 2.19 0.62 2.19  ;
        POLYGON 10.015 1.765 17.92 1.765 17.92 2.19 10.015 2.19  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.4624 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 2.42 8.79 2.42 8.79 1.445 1.365 1.445 1.365 0.675 1.625 0.675 1.625 0.865 3.605 0.865 3.605 0.675 3.835 0.675 3.835 0.865 5.845 0.865 5.845 0.675 6.075 0.675 6.075 0.865 8.085 0.865 8.085 0.675 8.315 0.675 8.315 0.865 10.325 0.865 10.325 0.675 10.555 0.675 10.555 0.865 12.565 0.865 12.565 0.675 12.795 0.675 12.795 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 1.445 9.69 1.445 9.69 2.42 17.175 2.42 17.175 3.39 16.945 3.39 16.945 3 14.935 3 14.935 3.39 14.705 3.39 14.705 3 12.695 3 12.695 3.39 12.465 3.39 12.465 3 10.455 3 10.455 3.39 10.225 3.39 10.225 3 8.31 3 8.31 3.39 8.08 3.39 8.08 3 5.975 3 5.975 3.39 5.745 3.39 5.745 3 3.735 3 3.735 3.39 3.505 3.39 3.505 3 1.595 3 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.68 0.475 2.68 0.475 3.62 2.385 3.62 2.385 3.23 2.615 3.23 2.615 3.62 4.625 3.62 4.625 3.23 4.855 3.23 4.855 3.62 6.865 3.62 6.865 3.23 7.095 3.23 7.095 3.62 9.105 3.62 9.105 3.23 9.335 3.23 9.335 3.62 11.345 3.62 11.345 3.23 11.575 3.23 11.575 3.62 13.585 3.62 13.585 3.23 13.815 3.23 13.815 3.62 15.825 3.62 15.825 3.23 16.055 3.23 16.055 3.62 18.065 3.62 18.065 2.68 18.295 2.68 18.295 3.62 19.04 3.62 19.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.395 0.3 18.395 1.015 18.165 1.015 18.165 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.73 0.3 11.73 0.635 11.39 0.635 11.39 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_16
