# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.85 1.45 2.87 1.45 2.87 1.795 3.52 1.795 4.27 1.795 4.27 1.265 4.565 1.265 4.565 2.095 3.52 2.095 2.595 2.095 2.595 1.68 1.85 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.915 1.8 1.61 1.8 1.61 1.91 2.315 1.91 2.315 2.325 3.52 2.325 4.83 2.325 4.83 1.8 6.225 1.8 6.225 2.12 5.105 2.12 5.105 2.68 3.52 2.68 3.375 2.68 3.375 2.555 2.035 2.555 2.035 2.14 0.915 2.14  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.195 2.36 9.08 2.36 9.315 2.36 9.315 1.56 8.195 1.56 8.195 0.61 8.545 0.61 8.545 1.24 9.6 1.24 9.6 2.68 9.08 2.68 8.56 2.68 8.56 3.38 8.195 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.455 3.62 0.455 2.83 0.685 2.83 0.685 3.62 2.72 3.62 2.72 2.79 3.06 2.79 3.06 3.62 3.52 3.62 6.32 3.62 6.32 2.815 6.66 2.815 6.66 3.62 7.295 3.62 7.295 2.53 7.525 2.53 7.525 3.62 9.08 3.62 9.335 3.62 9.335 2.94 9.565 2.94 9.565 3.62 10.08 3.62 10.08 4.22 9.08 4.22 3.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.665 0.3 9.665 0.99 9.435 0.99 9.435 0.3 7.425 0.3 7.425 0.99 7.195 0.99 7.195 0.3 2.96 0.3 2.96 0.76 2.62 0.76 2.62 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.4 0.53 0.74 0.53 0.74 0.99 3.52 0.99 3.52 1.555 3.18 1.555 3.18 1.22 0.68 1.22 0.68 2.37 1.705 2.37 1.705 3.35 1.475 3.35 1.475 2.6 0.4 2.6  ;
        POLYGON 3.65 0.53 6.77 0.53 6.77 0.76 3.65 0.76  ;
        POLYGON 3.6 2.99 5.4 2.99 5.4 2.35 6.54 2.35 6.54 1.22 5.07 1.22 5.07 0.99 6.77 0.99 6.77 1.82 9.08 1.82 9.08 2.095 6.77 2.095 6.77 2.58 5.63 2.58 5.63 3.22 3.6 3.22  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_2
