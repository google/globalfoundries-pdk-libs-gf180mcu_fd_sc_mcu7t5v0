* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
M_i_2_1 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 ZN B VDD VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_5_0 VDD B ZN VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_4_1 net_1_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_1 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_0 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 VDD A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS
