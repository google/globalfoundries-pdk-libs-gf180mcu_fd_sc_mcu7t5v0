# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__hold 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.4512 ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.565 0.475 0.565 0.475 1.155 3.95 1.155 3.95 1.56 0.575 1.56 0.575 2.895 0.245 2.895  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 3.225 3.62 3.225 2.535 3.455 2.535 3.455 3.62 4.575 3.62 5.04 3.62 5.04 4.22 4.575 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 3.455 0.3 3.455 0.925 3.225 0.925 3.225 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.45 1.885 4.345 1.885 4.345 0.575 4.575 0.575 4.575 3.18 4.245 3.18 4.245 2.185 2.45 2.185  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__hold
