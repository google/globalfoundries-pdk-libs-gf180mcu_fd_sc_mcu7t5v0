# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.955 1.825 4.39 1.825 4.39 2.095 2.955 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.77 2.385 1.77 2.385 1.36 4.895 1.36 4.895 1.77 5.65 1.77 5.65 2.15 4.625 2.15 4.625 1.59 2.71 1.59 2.71 2.095 1.935 2.095  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.39 1.58 1.39 1.58 2.38 6.25 2.38 6.25 1.73 6.63 1.73 6.63 2.655 1.305 2.655 1.305 1.665 0.705 1.665  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6492 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 0.53 0.53 0.53 0.53 0.885 1.89 0.885 1.89 0.53 3.31 0.53 3.31 0.885 4.13 0.885 4.13 0.53 5.55 0.53 5.55 0.885 6.905 0.885 6.905 0.53 7.25 0.53 7.25 1.115 0.42 1.115 0.42 2.02 1.055 2.02 1.055 2.94 3.84 2.94 3.84 3.235 0.825 3.235 0.825 2.25 0.145 2.25  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.59 0.575 2.59 0.575 3.62 6.865 3.62 6.865 2.63 7.095 2.63 7.095 3.62 7.84 3.62 7.84 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 6.14 0.3 6.14 0.655 5.78 0.655 5.78 0.3 3.9 0.3 3.9 0.655 3.54 0.655 3.54 0.3 1.66 0.3 1.66 0.655 1.3 0.655 1.3 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_2
