# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.6 2.13 0.6 2.13 1.79 2.855 1.79 2.855 2.13 1.825 2.13  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.18 1.01 1.18 1.01 3.32 0.705 3.32  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8306 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.6 1.595 0.6 1.595 2.36 2.665 2.36 2.665 3.38 2.385 3.38 2.385 2.68 1.24 2.68  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 3.36 3.62 3.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 2.715 0.3 2.715 1.09 2.485 1.09 2.485 0.3 0.475 0.3 0.475 0.945 0.245 0.945 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_1
