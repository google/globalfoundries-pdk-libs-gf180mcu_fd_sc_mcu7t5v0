# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.615 1.77 3.47 1.77 3.47 2.15 1.615 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.64 1.795 17.07 1.795 17.07 2.15 14.64 2.15  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.694 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.89 1.62 8.415 1.62 12.34 1.62 12.34 1.2 13.21 1.2 13.54 1.2 13.54 0.55 13.91 0.55 13.91 1.85 13.21 1.85 8.415 1.85 3.89 1.85  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 0.79 17.83 0.79 17.83 3.37 17.45 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.847 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.61 0.575 0.61 0.575 3.37 0.14 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.04 1.595 3.04 1.595 3.62 4.71 3.62 6.79 3.62 6.79 3.005 7.13 3.005 7.13 3.62 8.37 3.62 9.105 3.62 9.105 2.705 9.335 2.705 9.335 3.62 11.31 3.62 11.31 3.005 11.65 3.005 11.65 3.62 13.43 3.62 16.445 3.62 16.445 2.48 16.675 2.48 16.675 3.62 17.2 3.62 18.48 3.62 18.48 4.22 17.2 4.22 13.43 4.22 8.37 4.22 4.71 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.675 0.3 16.675 0.765 16.445 0.765 16.445 0.3 11.65 0.3 11.65 0.915 11.31 0.915 11.31 0.3 9.59 0.3 9.59 1.09 9.25 1.09 9.25 0.3 7.13 0.3 7.13 0.915 6.79 0.915 6.79 0.3 1.595 0.3 1.595 0.87 1.365 0.87 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.155 2.56 4.71 2.56 4.71 2.79 0.925 2.79 0.925 1.16 4.385 1.16 4.385 0.81 4.615 0.81 4.615 1.39 1.155 1.39  ;
        POLYGON 5.55 2.545 8.37 2.545 8.37 2.845 8.03 2.845 8.03 2.775 5.89 2.775 5.89 2.845 5.55 2.845  ;
        POLYGON 5.505 0.81 5.735 0.81 5.735 1.145 8.185 1.145 8.185 0.81 8.415 0.81 8.415 1.375 5.505 1.375  ;
        POLYGON 10.025 0.77 10.255 0.77 10.255 1.145 11.88 1.145 11.88 0.68 13.21 0.68 13.21 0.915 12.11 0.915 12.11 1.375 10.025 1.375  ;
        POLYGON 10.07 2.545 13.43 2.545 13.43 2.775 10.07 2.775  ;
        POLYGON 5.01 2.08 14.17 2.08 14.17 0.75 14.495 0.75 14.495 1.335 17.2 1.335 17.2 1.565 14.4 1.565 14.4 2.765 14.165 2.765 14.165 2.315 5.01 2.315  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_1
