# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.8 6.42 1.8 6.42 2.12 0.6 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.21 3.465 1.21 3.465 1.325 7.065 1.325 7.065 1.805 8.35 1.805 8.35 2.12 6.835 2.12 6.835 1.57 0.6 1.57  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.624 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.295 1.79 12.79 1.79 12.79 2.15 9.295 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.8792 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.41 2.38 8.58 2.38 8.58 1.475 7.765 1.475 7.765 1.095 3.87 1.095 3.87 0.825 2.37 0.825 2.37 0.595 4.1 0.595 4.1 0.865 7.995 0.865 7.995 1.245 9.605 1.245 9.605 0.655 9.835 0.655 9.835 1.245 11.845 1.245 11.845 0.655 12.075 0.655 12.075 1.56 8.87 1.56 8.87 2.765 1.41 2.765  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 9.85 3.62 9.85 3.04 10.19 3.04 10.19 3.62 11.89 3.62 11.89 3.04 12.23 3.04 12.23 3.62 13.25 3.62 13.44 3.62 13.44 4.22 13.25 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 13.195 0.3 13.195 1.215 12.965 1.215 12.965 0.3 11.01 0.3 11.01 1.015 10.67 1.015 10.67 0.3 8.59 0.3 8.59 0.98 8.25 0.98 8.25 0.3 4.67 0.3 4.67 0.635 4.33 0.635 4.33 0.3 0.695 0.3 0.695 0.69 0.465 0.69 0.465 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.445 2.54 0.675 2.54 0.675 3.16 9.235 3.16 9.235 2.53 13.25 2.53 13.25 3.38 12.91 3.38 12.91 2.76 11.21 2.76 11.21 3.38 10.87 3.38 10.87 2.76 9.565 2.76 9.565 3.39 0.445 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_4
