# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.66 1.085 1.02 1.085 1.02 2.87 0.66 2.87  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.78 1.58 2.26 1.58 2.26 3.28 1.78 3.28  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.9 1.58 3.38 1.58 3.38 3.28 2.9 3.28  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.02 1.58 4.5 1.58 4.5 3.28 4.02 3.28  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.07 0.63 6.575 0.63 6.575 3.38 6.07 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 5.085 3.62 5.085 2.53 5.315 2.53 5.315 3.62 5.765 3.62 6.72 3.62 6.72 4.22 5.765 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 5.315 0.3 5.315 0.855 5.085 0.855 5.085 0.3 2.95 0.3 2.95 0.76 2.61 0.76 2.61 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.28 3.12 1.3 3.12 1.3 1.095 1.49 1.095 1.49 0.53 1.83 0.53 1.83 1.095 3.73 1.095 3.73 0.53 4.07 0.53 4.07 1.095 5.765 1.095 5.765 2.27 5.515 2.27 5.515 1.33 1.53 1.33 1.53 3.35 0.28 3.35  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_1
