# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.694 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.74 2.855 1.74 2.855 2.12 0.65 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.754 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 3.46 2.36 3.46 1.505 1.365 1.505 1.365 0.7 1.595 0.7 1.595 1.27 3.45 1.27 3.45 0.65 3.835 0.65 3.835 3.38 3.45 3.38 3.45 2.735 1.495 2.735 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.55 0.475 2.55 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_3
