# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.715 1.74 3.78 1.74 3.78 2.35 7.38 2.35 7.38 2.205 7.77 2.205 7.77 2.71 3.435 2.71 3.435 2.15 2.715 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.21 4.39 1.21 4.39 1.72 5.62 1.72 5.62 2.12 4.01 2.12  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1771 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 0.55 1.615 0.55 1.615 3.37 1.21 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9308 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.49 2.25 10.79 2.25 11.31 2.25 11.31 1.56 10.49 1.56 10.49 0.55 11.11 0.55 11.11 1.22 11.65 1.22 11.65 2.48 11.11 2.48 11.11 3.37 10.79 3.37 10.49 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.315 3.62 0.315 2.48 0.545 2.48 0.545 3.62 2.4 3.62 2.4 3.215 2.74 3.215 2.74 3.62 4.49 3.62 4.49 3.215 4.83 3.215 4.83 3.62 5.43 3.62 5.43 3.215 5.77 3.215 5.77 3.62 9.37 3.62 9.37 2.685 9.71 2.685 9.71 3.62 10.79 3.62 11.51 3.62 11.51 2.71 11.85 2.71 11.85 3.62 12.32 3.62 12.32 4.22 10.79 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.895 0.3 11.895 0.78 11.665 0.78 11.665 0.3 9.655 0.3 9.655 0.78 9.425 0.78 9.425 0.3 2.735 0.3 2.735 0.94 2.505 0.94 2.505 0.3 0.495 0.3 0.495 0.985 0.265 0.985 0.265 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.33 0.53 8.35 0.53 8.35 0.76 5.33 0.76  ;
        POLYGON 2.015 1.18 3.125 1.18 3.125 0.53 4.895 0.53 4.895 1.19 6.325 1.19 6.325 1.745 8.79 1.745 8.79 1.975 6.095 1.975 6.095 1.42 4.665 1.42 4.665 0.76 3.355 0.76 3.355 1.41 2.245 1.41 2.245 2.755 3.205 2.755 3.205 2.94 3.81 2.94 3.81 3.17 2.975 3.17 2.975 2.985 2.015 2.985  ;
        POLYGON 8.01 2.205 9.17 2.205 9.17 1.515 6.67 1.515 6.67 0.99 7.01 0.99 7.01 1.285 9.4 1.285 9.4 1.79 10.79 1.79 10.79 2.02 9.4 2.02 9.4 2.435 8.35 2.435 8.35 3.37 8.01 3.37  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_2
