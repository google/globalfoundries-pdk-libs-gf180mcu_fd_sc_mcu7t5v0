# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.738 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.37 1.74 8.31 1.74 8.31 2.15 0.37 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.0688 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.505 2.42 17.16 2.42 17.985 2.42 17.985 1.535 10.505 1.535 10.505 0.69 10.735 0.69 10.735 1.215 12.745 1.215 12.745 0.69 12.975 0.69 12.975 1.215 14.985 1.215 14.985 0.69 15.215 0.69 15.215 1.215 17.225 1.215 17.225 0.69 17.455 0.69 17.455 1.215 19.465 1.215 19.465 0.69 19.695 0.69 19.695 1.215 21.705 1.215 21.705 0.69 21.935 0.69 21.935 1.215 23.945 1.215 23.945 0.69 24.175 0.69 24.175 1.215 26.185 1.215 26.185 0.69 26.415 0.69 26.415 1.535 18.885 1.535 18.885 2.42 26.315 2.42 26.315 3.39 26.085 3.39 26.085 3 24.075 3 24.075 3.39 23.845 3.39 23.845 3 21.835 3 21.835 3.39 21.605 3.39 21.605 3 19.595 3 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.16 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 12.875 3 12.875 3.39 12.645 3.39 12.645 3 10.735 3 10.735 3.39 10.505 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.865 3.62 6.865 3.05 7.095 3.05 7.095 3.62 9.385 3.62 9.385 3.19 9.615 3.19 9.615 3.62 11.525 3.62 11.525 3.23 11.755 3.23 11.755 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 17.16 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.485 3.62 20.485 3.23 20.715 3.23 20.715 3.62 22.725 3.62 22.725 3.23 22.955 3.23 22.955 3.62 24.965 3.62 24.965 3.23 25.195 3.23 25.195 3.62 27.16 3.62 27.205 3.62 27.205 2.76 27.435 2.76 27.435 3.62 28 3.62 28 4.22 27.16 4.22 17.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 28 -0.3 28 0.3 27.59 0.3 27.59 0.985 27.25 0.985 27.25 0.3 25.35 0.3 25.35 0.985 25.01 0.985 25.01 0.3 23.11 0.3 23.11 0.985 22.77 0.985 22.77 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.96 9.33 0.96 9.33 0.3 7.25 0.3 7.25 1.04 6.91 1.04 6.91 0.3 5.01 0.3 5.01 1.04 4.67 1.04 4.67 0.3 2.77 0.3 2.77 1.04 2.43 1.04 2.43 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 8.62 2.53 8.62 1.5 1.365 1.5 1.365 0.74 1.595 0.74 1.595 1.27 3.605 1.27 3.605 0.74 3.835 0.74 3.835 1.27 5.845 1.27 5.845 0.74 6.075 0.74 6.075 1.27 8.085 1.27 8.085 0.74 8.315 0.74 8.315 1.27 8.85 1.27 8.85 1.765 17.16 1.765 17.16 2.065 8.85 2.065 8.85 2.76 8.215 2.76 8.215 3.39 7.985 3.39 7.985 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.495 2.76 1.495 3.39 1.265 3.39  ;
        POLYGON 19.74 1.765 27.16 1.765 27.16 2.065 19.74 2.065  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
