* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
M_MN2_12 VSS int04 Z VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN2 VSS int04 Z VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN4 net_1 I1 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN8 int04 S net_1 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN7 net_3 sel1_n int04 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN3 VSS I0 net_3 VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MN1 sel1_n S VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_MP5_6 VDD int04 Z VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP5 VDD int04 Z VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP4 net_0 I1 VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP8 int04 sel1_n net_0 VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP7 net_2 S int04 VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP3 VDD I0 net_2 VNW pmos_5p0 W=1.22e-06 L=5e-07
M_MP1 sel1_n S VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
