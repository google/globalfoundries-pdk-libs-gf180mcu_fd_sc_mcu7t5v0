# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.77 1.56 1.77 1.56 2.19 1 2.19 1 3 0.66 3  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.015 1.21 2.13 1.21 2.13 2.41 1.79 2.41 1.79 1.54 1.015 1.54  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 1.21 3.43 1.21 3.43 1.57 2.7 1.57 2.7 2.41 2.36 2.41  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.215 1.8 4.78 1.8 4.78 2.12 3.215 2.12  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.66 0.61 6.03 0.61 6.03 3.35 5.66 3.35  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.25 3.62 0.25 3.285 0.59 3.285 0.59 3.62 2.29 3.62 2.29 3.285 2.63 3.285 2.63 3.62 4.55 3.62 4.55 3.285 4.89 3.285 4.89 3.62 5.385 3.62 6.16 3.62 6.16 4.22 5.385 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 4.845 0.3 4.845 1.035 4.505 1.035 4.505 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.27 2.825 5.155 2.825 5.155 1.505 3.77 1.505 3.77 0.76 0.535 0.76 0.535 1.09 0.305 1.09 0.305 0.53 4 0.53 4 1.265 5.385 1.265 5.385 3.055 3.65 3.055 3.65 3.39 3.31 3.39 3.31 3.055 1.61 3.055 1.61 3.39 1.27 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_1
