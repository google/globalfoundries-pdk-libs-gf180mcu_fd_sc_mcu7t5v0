# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.306 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.41 1.76 3.015 1.76 3.015 2.12 0.41 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2024 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 2.36 3.41 2.36 3.41 1.525 1.365 1.525 1.365 0.53 1.595 0.53 1.595 1.29 3.41 1.29 3.41 0.53 3.835 0.53 3.835 3.39 3.41 3.39 3.41 2.68 1.595 2.68 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.485 3.62 2.485 2.985 2.715 2.985 2.715 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.055 2.485 1.055 2.485 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_3
