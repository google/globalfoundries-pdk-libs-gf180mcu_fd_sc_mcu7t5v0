# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.2 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.775 1.63 1.775 1.63 2.185 0.545 2.185  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.09 1.8 7.275 1.8 7.275 2.12 5.09 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9152 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.46 2.54 10.37 2.54 10.49 2.54 10.74 2.54 10.74 1.135 8.34 1.135 8.34 0.865 11.07 0.865 11.07 2.77 10.84 2.77 10.84 3.39 10.5 3.39 10.5 2.77 10.49 2.77 10.37 2.77 8.8 2.77 8.8 3.39 8.46 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.22 3.62 5.22 3.285 5.56 3.285 5.56 3.62 7.26 3.62 7.26 3.285 7.6 3.285 7.6 3.62 9.48 3.62 9.48 3.285 9.82 3.285 9.82 3.62 10.37 3.62 10.49 3.62 11.2 3.62 11.2 4.22 10.49 4.22 10.37 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.2 -0.3 11.2 0.3 9.89 0.3 9.89 0.635 9.55 0.635 9.55 0.3 7.56 0.3 7.56 0.635 7.22 0.635 7.22 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.925 2.78 1.925 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.155 1.095 2.155 2.235 3.65 2.235 3.65 2.52 2.155 2.52 2.155 3.01 0.42 3.01  ;
        POLYGON 2.87 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.575 7.625 2.575 7.625 1.965 10.37 1.965 10.37 2.195 7.855 2.195 7.855 2.805 6.58 2.805 6.58 3.39 6.24 3.39 6.24 2.805 4.825 2.805 4.825 3.39 2.87 3.39  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 5.92 0.705 5.92 0.585 6.37 0.585 6.37 0.865 8.015 0.865 8.015 1.365 10.49 1.365 10.49 1.595 7.785 1.595 7.785 1.095 5.92 1.095 5.92 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_3
