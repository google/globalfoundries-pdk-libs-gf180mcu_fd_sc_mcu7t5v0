# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4565 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.85 1.65 3.96 1.65 3.96 2.15 2.85 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.177 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.715 1.785 18.115 1.785 18.115 2.13 16.715 2.13  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.565 1.67 15.955 1.67 15.955 2.225 14.565 2.225  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 0.6 1.07 0.6 1.07 2.15 0.705 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1112 ;
    PORT
      LAYER METAL1 ;
        POLYGON 21.045 2.125 22.89 2.125 23.14 2.125 23.14 1.315 21.045 1.315 21.045 0.655 21.275 0.655 21.275 1.085 23.14 1.085 23.14 0.6 24.005 0.6 24.005 2.28 23.42 2.28 23.42 3.38 23.06 3.38 23.06 2.36 22.89 2.36 21.335 2.36 21.335 3.38 21.045 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.205 3.62 1.205 2.93 1.555 2.93 1.555 3.62 2.035 3.62 3.01 3.62 3.01 3.005 3.35 3.005 3.35 3.62 4.995 3.62 7.53 3.62 7.53 3.445 7.87 3.445 7.87 3.62 10.73 3.62 10.73 3.445 11.07 3.445 11.07 3.62 12.75 3.62 15.125 3.62 15.125 2.93 15.465 2.93 15.465 3.62 17.27 3.62 17.27 2.93 17.61 2.93 17.61 3.62 19.035 3.62 19.365 3.62 19.365 2.73 19.595 2.73 19.595 3.62 20.085 3.62 20.085 2.53 20.315 2.53 20.315 3.62 22.07 3.62 22.07 2.62 22.41 2.62 22.41 3.62 22.89 3.62 24.165 3.62 24.165 2.53 24.395 2.53 24.395 3.62 25.2 3.62 25.2 4.22 22.89 4.22 19.035 4.22 12.75 4.22 4.995 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 24.635 0.3 24.635 0.905 24.405 0.905 24.405 0.3 22.395 0.3 22.395 0.765 22.165 0.765 22.165 0.3 20.155 0.3 20.155 0.905 19.925 0.905 19.925 0.3 17.51 0.3 17.51 1.075 17.17 1.075 17.17 0.3 9.19 0.3 9.19 0.915 8.85 0.915 8.85 0.3 3.85 0.3 3.85 1.15 3.51 1.15 3.51 0.3 1.595 0.3 1.595 1.16 1.365 1.16 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.81 0.475 0.81 0.475 2.38 1.805 2.38 1.805 1.28 2.035 1.28 2.035 2.7 0.475 2.7 0.475 3.225 0.245 3.225  ;
        POLYGON 4.305 0.865 4.915 0.865 4.915 1.205 4.535 1.205 4.535 2.93 4.305 2.93  ;
        POLYGON 2.515 2.49 3.88 2.49 3.88 3.16 4.765 3.16 4.765 1.895 4.995 1.895 4.995 3.39 3.65 3.39 3.65 2.725 2.515 2.725 2.515 3.225 2.285 3.225 2.285 0.765 2.715 0.765 2.715 1.105 2.515 1.105  ;
        POLYGON 6.29 2.525 9.11 2.525 9.11 2.93 8.77 2.93 8.77 2.755 6.63 2.755 6.63 2.885 6.29 2.885  ;
        POLYGON 5.325 2.04 5.805 2.04 5.805 0.865 6.035 0.865 6.035 2.065 10.36 2.065 10.36 2.295 5.555 2.295 5.555 2.94 5.325 2.94  ;
        POLYGON 9.49 2.525 11.28 2.525 11.28 1.835 7.03 1.835 7.03 1.605 11.17 1.605 11.17 0.99 11.51 0.99 11.51 2.525 12.31 2.525 12.31 2.835 11.97 2.835 11.97 2.755 9.83 2.755 9.83 2.93 9.49 2.93  ;
        POLYGON 5.78 3.16 7.07 3.16 7.07 2.985 8.41 2.985 8.41 3.16 10.245 3.16 10.245 2.985 11.53 2.985 11.53 3.065 12.75 3.065 12.75 3.295 11.3 3.295 11.3 3.215 10.48 3.215 10.48 3.39 8.18 3.39 8.18 3.215 7.3 3.215 7.3 3.39 5.78 3.39  ;
        POLYGON 6.265 1.145 10.65 1.145 10.65 0.53 13.125 0.53 13.125 1.6 13.735 1.6 13.735 2.43 13.505 2.43 13.505 1.83 12.895 1.83 12.895 0.76 12 0.76 12 1.735 11.745 1.735 11.745 0.76 10.88 0.76 10.88 1.375 6.495 1.375 6.495 1.685 6.265 1.685  ;
        POLYGON 13.41 0.99 14.065 0.99 14.065 0.845 16.415 0.845 16.415 2.465 16.535 2.465 16.535 2.805 16.185 2.805 16.185 1.075 14.295 1.075 14.295 2.89 14.065 2.89 14.065 1.22 13.41 1.22  ;
        POLYGON 12.29 0.99 12.63 0.99 12.63 2.06 13.275 2.06 13.275 3.12 14.585 3.12 14.585 2.465 15.925 2.465 15.925 3.09 16.805 3.09 16.805 2.465 18.115 2.465 18.115 3.035 18.805 3.035 18.805 2.005 19.035 2.005 19.035 3.27 17.885 3.27 17.885 2.7 17.035 2.7 17.035 3.325 15.695 3.325 15.695 2.7 14.815 2.7 14.815 3.355 13.045 3.355 13.045 2.295 12.4 2.295 12.4 1.22 12.29 1.22  ;
        POLYGON 16.645 1.325 19.205 1.325 19.205 0.79 19.435 0.79 19.435 1.325 20.595 1.325 20.595 1.555 22.89 1.555 22.89 1.785 20.305 1.785 20.305 1.555 18.575 1.555 18.575 2.805 18.345 2.805 18.345 1.555 16.645 1.555  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
