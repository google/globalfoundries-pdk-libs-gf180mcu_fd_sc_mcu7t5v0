# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.816 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.71 8.185 1.71 8.185 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.4624 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.325 2.23 16.51 2.23 17.75 2.23 17.75 1.51 10.325 1.51 10.325 0.675 10.585 0.675 10.585 0.93 12.565 0.93 12.565 0.675 12.795 0.675 12.795 0.93 14.805 0.93 14.805 0.675 15.035 0.675 15.035 0.93 17.045 0.93 17.045 0.675 17.275 0.675 17.275 0.93 19.285 0.93 19.285 0.675 19.515 0.675 19.515 0.93 21.525 0.93 21.525 0.675 21.755 0.675 21.755 0.93 23.765 0.93 23.765 0.675 23.995 0.675 23.995 0.93 26.005 0.93 26.005 0.675 26.235 0.675 26.235 1.51 18.65 1.51 18.65 2.23 26.135 2.23 26.135 3.38 25.905 3.38 25.905 2.81 23.895 2.81 23.895 3.38 23.665 3.38 23.665 2.81 21.655 2.81 21.655 3.38 21.425 3.38 21.425 2.81 19.415 2.81 19.415 3.38 19.185 3.38 19.185 2.81 17.175 2.81 17.175 3.38 16.945 3.38 16.945 2.81 16.51 2.81 14.935 2.81 14.935 3.38 14.705 3.38 14.705 2.81 12.695 2.81 12.695 3.38 12.465 3.38 12.465 2.81 10.555 2.81 10.555 3.38 10.325 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 3 7.095 3 7.095 3.62 9.105 3.62 9.105 2.53 9.335 2.53 9.335 3.62 11.345 3.62 11.345 3.04 11.575 3.04 11.575 3.62 13.585 3.62 13.585 3.04 13.815 3.04 13.815 3.62 15.825 3.62 15.825 3.04 16.055 3.04 16.055 3.62 16.51 3.62 18.065 3.62 18.065 3.04 18.295 3.04 18.295 3.62 20.305 3.62 20.305 3.04 20.535 3.04 20.535 3.62 22.545 3.62 22.545 3.04 22.775 3.04 22.775 3.62 24.785 3.62 24.785 3.04 25.015 3.04 25.015 3.62 26.98 3.62 27.025 3.62 27.025 2.53 27.255 2.53 27.255 3.62 28 3.62 28 4.22 26.98 4.22 16.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 28 -0.3 28 0.3 27.41 0.3 27.41 0.765 27.07 0.765 27.07 0.3 25.17 0.3 25.17 0.7 24.83 0.7 24.83 0.3 22.93 0.3 22.93 0.7 22.59 0.7 22.59 0.3 20.69 0.3 20.69 0.7 20.35 0.7 20.35 0.3 18.45 0.3 18.45 0.7 18.11 0.7 18.11 0.3 16.21 0.3 16.21 0.7 15.87 0.7 15.87 0.3 13.97 0.3 13.97 0.7 13.63 0.7 13.63 0.3 11.73 0.3 11.73 0.7 11.39 0.7 11.39 0.3 9.49 0.3 9.49 0.765 9.15 0.765 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 8.535 2.53 8.535 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 5.845 1.015 5.845 0.675 6.075 0.675 6.075 1.015 8.085 1.015 8.085 0.675 8.315 0.675 8.315 1.015 8.77 1.015 8.77 1.74 16.51 1.74 16.51 1.97 8.77 1.97 8.77 2.76 8.215 2.76 8.215 3.38 7.985 3.38 7.985 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 19.56 1.74 26.98 1.74 26.98 1.97 19.56 1.97  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_16
