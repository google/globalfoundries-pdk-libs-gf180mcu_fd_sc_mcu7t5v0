# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.91 1.575 3.25 1.575 3.25 3.39 2.91 3.39  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 1.575 2.13 1.575 2.13 3.39 1.79 3.39  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.49 1.76 1.56 1.76 1.56 3.39 1.22 3.39 1.22 2.19 0.49 2.19  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9832 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.31 0.695 1.65 0.695 1.65 1.05 3.55 1.05 3.55 0.695 3.89 0.695 3.89 3.39 3.49 3.39 3.49 1.285 1.31 1.285  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.77 0.3 2.77 0.82 2.43 0.82 2.43 0.3 0.53 0.3 0.53 0.82 0.19 0.82 0.19 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_1
