* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addf_1 A B CI CO S VDD VNW VPW VSS
M_M51 VSS net9 S VPW nmos_5p0 W=7.1e-07 L=6e-07
M_M46 net9 CI net47 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M45 net42 CI VSS VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M34 CO net7 VSS VPW nmos_5p0 W=8.15e-07 L=6e-07
M_M33 VDD net9 S VNW pmos_5p0 W=1.215e-06 L=5e-07
M_M28 net9 CI net29 VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M24 net9 net7 net3 VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M25 net3 A VDD VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M26 VDD B net3 VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M27 net3 CI VDD VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M21 net7 CI net1 VNW pmos_5p0 W=7e-07 L=5e-07
M_M20 net19 B net7 VNW pmos_5p0 W=7e-07 L=5e-07
M_M18 VDD A net19 VNW pmos_5p0 W=7e-07 L=5e-07
M_M17 CO net7 VDD VNW pmos_5p0 W=1.215e-06 L=5e-07
M_M48 net47 B net49 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M41 net9 net7 net42 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M43 net42 A VSS VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M44 VSS B net42 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M38 net7 CI net5 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M37 net36 B net7 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M35 VSS A net36 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M30 net29 B net31 VNW pmos_5p0 W=6.6e-07 L=5e-07
M_M23 VDD B net1 VNW pmos_5p0 W=7e-07 L=5e-07
M_M22 net1 A VDD VNW pmos_5p0 W=7e-07 L=5e-07
M_M50 net49 A VSS VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M40 VSS B net5 VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M39 net5 A VSS VPW nmos_5p0 W=3.8e-07 L=6e-07
M_M32 net31 A VDD VNW pmos_5p0 W=6.6e-07 L=5e-07
.ENDS
