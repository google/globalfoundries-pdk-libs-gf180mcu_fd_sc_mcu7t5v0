# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.555 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.765 6.07 1.765 6.07 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.036 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.265 2.495 13.09 2.495 13.83 2.495 13.83 1.535 8.265 1.535 8.265 0.69 8.495 0.69 8.495 1.215 10.505 1.215 10.505 0.69 10.735 0.69 10.735 1.215 12.745 1.215 12.745 0.69 12.975 0.69 12.975 1.215 14.985 1.215 14.985 0.69 15.215 0.69 15.215 1.215 17.225 1.215 17.225 0.69 17.455 0.69 17.455 1.215 19.465 1.215 19.465 0.69 19.695 0.69 19.695 1.535 14.73 1.535 14.73 2.495 19.595 2.495 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 13.09 3 12.875 3 12.875 3.39 12.645 3.39 12.645 3 10.635 3 10.635 3.39 10.405 3.39 10.405 3 8.495 3 8.495 3.39 8.265 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 7.145 3.62 7.145 3.23 7.375 3.23 7.375 3.62 9.285 3.62 9.285 3.23 9.515 3.23 9.515 3.62 11.525 3.62 11.525 3.23 11.755 3.23 11.755 3.62 13.09 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.43 3.62 20.485 3.62 20.485 2.76 20.715 2.76 20.715 3.62 21.28 3.62 21.28 4.22 20.43 4.22 13.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.985 9.33 0.985 9.33 0.3 7.43 0.3 7.43 1.075 7.09 1.075 7.09 0.3 5.01 0.3 5.01 1.075 4.67 1.075 4.67 0.3 2.77 0.3 2.77 1.075 2.43 1.075 2.43 0.3 0.53 0.3 0.53 1.075 0.19 1.075 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 6.365 2.53 6.365 1.535 1.31 1.535 1.31 0.845 1.65 0.845 1.65 1.305 3.55 1.305 3.55 0.845 3.89 0.845 3.89 1.305 5.79 1.305 5.79 0.845 6.13 0.845 6.13 1.305 6.595 1.305 6.595 1.765 13.09 1.765 13.09 2.065 6.595 2.065 6.595 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.495 2.76 1.495 3.39 1.265 3.39  ;
        POLYGON 15.39 1.765 20.43 1.765 20.43 2.065 15.39 2.065  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
