# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.8 BY 3.92 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.679 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.11 1.535 10.74 1.535 10.74 1.21 11.235 1.21 12.755 1.21 12.755 1.59 11.235 1.59 10.97 1.59 10.97 1.765 10.11 1.765  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.8 2.75 1.8 2.75 3.37 2.34 3.37 2.34 2.12 1.865 2.12  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.8 1.59 1.8 1.59 2.12 0.29 2.12  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.118 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 2.4 14.97 2.4 15.22 2.4 15.22 1.08 14.555 1.08 14.555 0.6 15.58 0.6 15.58 2.74 15.02 2.74 15.02 3.38 14.97 3.38 14.66 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.29 3.62 0.29 2.535 0.63 2.535 0.63 3.62 2.77 3.62 6.28 3.62 6.28 2.505 6.51 2.505 6.51 3.62 9.69 3.62 9.69 2.92 9.92 2.92 9.92 3.62 11.635 3.62 11.635 2.57 11.865 2.57 11.865 3.62 13.645 3.62 13.645 2.815 13.985 2.815 13.985 3.62 14.97 3.62 15.87 3.62 15.87 2.53 16.1 2.53 16.1 3.62 16.8 3.62 16.8 4.22 14.97 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 16.8 -0.3 16.8 0.3 16.235 0.3 16.235 0.75 15.885 0.75 15.885 0.3 13.93 0.3 13.93 0.845 13.7 0.845 13.7 0.3 10.05 0.3 10.05 0.845 9.82 0.845 9.82 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 0.995 1.31 0.995 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.765 0.53 0.765 0.53 1.225 1.885 1.225 1.885 0.765 2.77 0.765 2.77 0.995 2.115 0.995 2.115 1.46 0.19 1.46  ;
        POLYGON 3.46 1.445 3.69 1.445 3.69 1.87 4.935 1.87 4.935 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 5.205 2.33 5.205 1.34 7.08 1.34 7.08 1.575 5.435 1.575 5.435 2.56 4.04 2.56 4.04 3.265 3.81 3.265 3.81 2.56 3 2.56 3 0.765 3.89 0.765 3.89 0.995 3.23 0.995  ;
        POLYGON 7.915 0.53 9.075 0.53 9.075 0.76 8.275 0.76 8.275 1.805 8.93 1.805 8.93 2.85 8.645 2.85 8.645 2.035 7.915 2.035  ;
        POLYGON 9.175 1.075 10.28 1.075 10.28 0.53 11.235 0.53 11.235 0.76 10.51 0.76 10.51 1.305 9.415 1.305 9.415 1.995 10.945 1.995 10.945 2.85 10.715 2.85 10.715 2.225 9.175 2.225  ;
        POLYGON 5.685 1.805 7.32 1.805 7.32 0.78 7.55 0.78 7.55 3.16 9.165 3.16 9.165 2.455 10.43 2.455 10.43 3.16 11.175 3.16 11.175 1.895 13.415 1.895 13.415 2.125 11.405 2.125 11.405 3.39 10.2 3.39 10.2 2.69 9.395 2.69 9.395 3.39 7.32 3.39 7.32 2.035 5.685 2.035  ;
        POLYGON 12.68 2.355 13.645 2.355 13.645 1.535 13.01 1.535 13.01 0.76 11.595 0.76 11.595 0.53 13.24 0.53 13.24 1.265 13.875 1.265 13.875 1.595 14.97 1.595 14.97 1.825 13.875 1.825 13.875 2.585 12.91 2.585 12.91 3.38 12.68 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_2
