# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.25 1.75 15.275 1.75 16.94 1.75 16.94 2.12 15.275 2.12 15.25 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.59 1.78 12.5 1.78 12.5 2.13 10.59 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.97 1.01 0.97 1.01 2.95 0.705 2.95  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.3 1.375 4.585 1.375 4.585 1.8 5.55 1.8 5.55 2.15 4.3 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.185 1.8 3.2 1.8 3.2 1.24 3.495 1.24 3.495 2.12 2.415 2.12 2.415 2.465 2.185 2.465  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.003 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.96 1.165 8.3 1.165 8.3 1.77 8.76 1.77 9.3 1.77 9.3 2.465 9.07 2.465 9.07 2.15 8.76 2.15 7.96 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.5104 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.65 0.6 6.38 0.6 6.38 2.855 5.99 2.855 5.99 1.57 5.65 1.57  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.685 0.475 2.685 0.475 3.62 1.65 3.62 4.845 3.62 4.845 2.845 5.185 2.845 5.185 3.62 7.27 3.62 8.76 3.62 11.67 3.62 11.67 2.845 12.015 2.845 12.015 3.62 14.1 3.62 15.955 3.62 15.955 2.815 16.295 2.815 16.295 3.62 17.46 3.62 17.92 3.62 17.92 4.22 17.46 4.22 14.1 4.22 8.76 4.22 7.27 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.34 0.3 16.34 1.145 16.11 1.145 16.11 0.3 11.86 0.3 11.86 1.145 11.63 1.145 11.63 0.3 5.08 0.3 5.08 1.16 4.85 1.16 4.85 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 3.025 1.26 3.025  ;
        POLYGON 3.725 0.78 4.07 0.78 4.07 2.87 3.725 2.87  ;
        POLYGON 6.86 2.665 7.27 2.665 7.27 3.005 6.86 3.005 6.86 3.39 5.52 3.39 5.52 2.615 4.53 2.615 4.53 3.33 2.635 3.33 2.635 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.77 0.845 2.77 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 2.975 2.74 2.975 3.1 4.3 3.1 4.3 2.38 5.75 2.38 5.75 3.155 6.63 3.155 6.63 0.79 7.27 0.79 7.27 1.13 6.86 1.13  ;
        POLYGON 7.09 1.46 7.5 1.46 7.5 0.53 8.76 0.53 8.76 1.145 8.53 1.145 8.53 0.76 7.73 0.76 7.73 2.72 8.755 2.72 8.755 2.95 7.5 2.95 7.5 1.82 7.09 1.82  ;
        POLYGON 10.35 2.575 10.84 2.575 10.84 2.925 10.11 2.925 10.11 0.795 10.84 0.795 10.84 1.145 10.35 1.145  ;
        POLYGON 12.75 0.78 12.98 0.78 12.98 2.925 12.75 2.925  ;
        POLYGON 9.65 0.78 9.88 0.78 9.88 3.16 11.125 3.16 11.125 2.38 12.495 2.38 12.495 3.16 13.77 3.16 13.77 0.78 14.1 0.78 14.1 3.39 12.265 3.39 12.265 2.615 11.355 2.615 11.355 3.39 9.65 3.39  ;
        POLYGON 14.33 0.85 15.275 0.85 15.275 1.08 14.56 1.08 14.56 2.815 15.19 2.815 15.19 3.045 14.33 3.045  ;
        POLYGON 14.79 1.685 15.02 1.685 15.02 2.355 17.23 2.355 17.23 0.78 17.46 0.78 17.46 3.14 17.125 3.14 17.125 2.585 14.79 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_1
