# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4985 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 0.65 1.22 0.65 1.22 1.63 1.59 1.63 1.59 2.19 0.705 2.19  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.33 0.575 2.955 0.575 2.955 3.38 2.485 3.38 2.485 1.6 2.33 1.6  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.53 3.62 1.53 3.13 1.87 3.13 1.87 3.62 2.255 3.62 3.36 3.62 3.36 4.22 2.255 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 1.815 0.3 1.815 0.865 1.585 0.865 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.8 0.475 0.8 0.475 2.58 1.97 2.58 1.97 1.83 2.255 1.83 2.255 2.815 0.63 2.815 0.63 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_1
