# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.394 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.81 1.21 13.865 1.21 13.865 1.45 14.255 1.45 14.255 2.195 14.025 2.195 14.025 1.68 13.57 1.68 13.57 1.59 11.81 1.59  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.845 1.77 2.73 1.77 2.73 3.37 2.32 3.37 2.32 2.15 1.845 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.27 1.77 1.57 1.77 1.57 2.15 0.27 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8118 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.3 0.63 17.035 0.63 17.035 3.27 16.3 3.27  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.3 3.62 6.3 2.79 6.53 2.79 6.53 3.62 8.79 3.62 9.11 3.62 9.11 2.47 9.34 2.47 9.34 3.62 9.91 3.62 12.8 3.62 12.8 2.46 13.03 2.46 13.03 3.62 13.63 3.62 15.345 3.62 15.345 2.425 15.685 2.425 15.685 3.62 16.07 3.62 17.36 3.62 17.36 4.22 16.07 4.22 13.63 4.22 9.91 4.22 8.79 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 15.91 0.3 15.91 1.095 15.68 1.095 15.68 0.3 15.245 0.3 15.245 0.76 14.905 0.76 14.905 0.3 13.005 0.3 13.005 0.76 12.665 0.76 12.665 0.3 9.445 0.3 9.445 1.075 9.105 1.075 9.105 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 1.06 1.31 1.06 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.845 0.53 0.845 0.53 1.29 1.885 1.29 1.885 0.845 2.77 0.845 2.77 1.075 2.115 1.075 2.115 1.52 0.19 1.52  ;
        POLYGON 3.46 1.42 3.69 1.42 3.69 1.87 7.32 1.87 7.32 0.78 7.55 0.78 7.55 2.9 7.32 2.9 7.32 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 7.04 2.33 7.04 3.16 8.56 3.16 8.56 1.82 8.79 1.82 8.79 3.39 6.81 3.39 6.81 2.56 4.04 2.56 4.04 3.125 3.81 3.125 3.81 2.56 3 2.56 3 0.845 3.89 0.845 3.89 1.075 3.23 1.075  ;
        POLYGON 8.04 0.78 8.27 0.78 8.27 1.34 9.91 1.34 9.91 1.575 8.27 1.575 8.27 2.9 8.04 2.9  ;
        POLYGON 11.09 2.26 12.01 2.26 12.01 2.93 11.78 2.93 11.78 2.495 10.86 2.495 10.86 0.53 11.975 0.53 11.975 0.76 11.09 0.76  ;
        POLYGON 10.18 0.78 10.51 0.78 10.51 3.16 12.34 3.16 12.34 1.91 13.63 1.91 13.63 2.14 12.57 2.14 12.57 3.39 10.18 3.39  ;
        POLYGON 13.785 0.53 14.57 0.53 14.57 0.99 14.79 0.99 14.79 1.79 16.07 1.79 16.07 2.13 14.79 2.13 14.79 3.18 14.56 3.18 14.56 1.22 14.34 1.22 14.34 0.76 13.785 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_1
