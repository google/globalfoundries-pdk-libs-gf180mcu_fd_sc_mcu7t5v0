# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.12 1.335 20.72 1.335 20.72 1.22 21.865 1.22 21.865 1.57 17.39 1.57 17.39 1.675 14.55 1.675 14.55 2.245 14.12 2.245  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.98 1.91 18.01 1.91 18.01 1.8 21.865 1.8 21.865 2.14 14.98 2.14  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.2 1.59 1.2 1.59 1.33 3.38 1.33 3.38 1.24 5.63 1.24 5.63 1.555 8.31 1.555 8.31 1.79 3.38 1.79 3.38 1.56 0.62 1.56  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.465 1.8 3.125 1.8 3.125 2.04 7.29 2.04 7.29 2.27 2.71 2.27 2.71 2.12 0.465 2.12  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.582 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.82 1.8 13.16 1.8 13.16 2.12 8.82 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.3055 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.73 2.05 0.73 2.05 0.87 2.85 0.87 2.85 0.545 6.11 0.545 6.11 1.095 8.555 1.095 8.555 0.765 8.785 0.765 8.785 1.095 11.11 1.095 11.11 0.53 11.45 0.53 11.45 1.095 13.53 1.095 13.53 0.53 13.87 0.53 13.87 0.875 16.24 0.875 16.24 0.545 18.69 0.545 18.69 0.87 20.24 0.87 20.24 0.545 22.04 0.545 22.04 0.775 20.47 0.775 20.47 1.105 18.46 1.105 18.46 0.78 16.47 0.78 16.47 1.105 13.88 1.105 13.88 2.68 21.05 2.68 21.05 2.91 13.53 2.91 13.53 1.56 8.905 1.56 8.905 1.325 5.88 1.325 5.88 0.78 3.08 0.78 3.08 1.1 1.82 1.1 1.82 0.96 0.19 0.96  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.24 3.62 0.24 2.53 0.58 2.53 0.58 3.62 2.335 3.62 2.335 3.04 2.565 3.04 2.565 3.62 4.375 3.62 4.375 3.04 4.605 3.04 4.605 3.62 6.415 3.62 6.415 3.04 6.645 3.04 6.645 3.62 8.455 3.62 8.455 3.04 8.685 3.04 8.685 3.62 21.975 3.62 22.4 3.62 22.4 4.22 21.975 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 19.99 0.3 19.99 0.64 19.65 0.64 19.65 0.3 15.91 0.3 15.91 0.64 15.57 0.64 15.57 0.3 12.515 0.3 12.515 0.795 12.285 0.795 12.285 0.3 10.275 0.3 10.275 0.795 10.045 0.795 10.045 0.3 6.7 0.3 6.7 0.795 6.36 0.795 6.36 0.3 2.62 0.3 2.62 0.64 2.28 0.64 2.28 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 2.53 12.56 2.53 12.56 2.76 7.72 2.76 7.72 3.38 7.38 3.38 7.38 2.76 5.68 2.76 5.68 3.38 5.34 3.38 5.34 2.76 3.64 2.76 3.64 3.38 3.3 3.38 3.3 2.76 1.6 2.76 1.6 3.38 1.26 3.38  ;
        POLYGON 9.11 3.16 21.745 3.16 21.745 2.5 21.975 2.5 21.975 3.39 9.11 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_4
