# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.795 5.14 1.795 5.14 2.215 3.41 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.739 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.465 1.795 6.63 1.795 6.63 2.2 5.465 2.2  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.11635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.76 0.615 21.18 0.615 21.18 3.39 20.76 3.39  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 2.775 3.62 5.25 3.62 5.25 3.18 5.59 3.18 5.59 3.62 7.57 3.62 7.57 3.35 7.91 3.35 7.91 3.62 10.015 3.62 12.93 3.62 12.93 2.995 13.27 2.995 13.27 3.62 16.245 3.62 17.71 3.62 17.71 2.8 18.05 2.8 18.05 3.62 18.63 3.62 19.785 3.62 19.785 2.46 20.015 2.46 20.015 3.62 20.515 3.62 21.875 3.62 21.875 2.46 22.105 2.46 22.105 3.62 22.4 3.62 22.4 4.22 20.515 4.22 18.63 4.22 16.245 4.22 10.015 4.22 2.775 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.155 0.3 22.155 0.95 21.925 0.95 21.925 0.3 19.915 0.3 19.915 0.95 19.685 0.95 19.685 0.3 18.075 0.3 18.075 0.725 17.845 0.725 17.845 0.3 13.32 0.3 13.32 1.085 12.98 1.085 12.98 0.3 8.01 0.3 8.01 1.045 7.78 1.045 7.78 0.3 5.635 0.3 5.635 1.075 5.295 1.075 5.295 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.385 2.545 2.385 2.545 1.625 2.775 1.625 2.775 2.615 0.475 2.615 0.475 3.015 0.245 3.015  ;
        POLYGON 6.585 2.43 6.86 2.43 6.86 1.275 6.75 1.275 6.75 0.99 7.09 0.99 7.09 2.43 8.37 2.43 8.37 1.875 8.6 1.875 8.6 2.66 6.815 2.66 6.815 2.86 6.585 2.86  ;
        POLYGON 3.03 2.705 6.105 2.705 6.105 3.09 7.09 3.09 7.09 2.89 8.6 2.89 8.6 3.12 9.785 3.12 9.785 2.69 10.015 2.69 10.015 3.35 8.37 3.35 8.37 3.12 7.32 3.12 7.32 3.32 5.875 3.32 5.875 2.935 3.03 2.935  ;
        POLYGON 3.27 0.845 4.655 0.845 4.655 1.305 6.035 1.305 6.035 0.53 7.55 0.53 7.55 1.305 8.375 1.305 8.375 0.53 10.07 0.53 10.07 1.14 9.84 1.14 9.84 0.76 8.605 0.76 8.605 1.535 7.32 1.535 7.32 0.76 6.265 0.76 6.265 1.535 4.425 1.535 4.425 1.075 3.27 1.075  ;
        POLYGON 10.855 1.47 10.96 1.47 10.96 0.8 11.19 0.8 11.19 1.47 13.965 1.47 13.965 1.7 11.085 1.7 11.085 2.87 10.855 2.87  ;
        POLYGON 12.2 2.07 14.285 2.07 14.285 0.8 14.555 0.8 14.555 2.87 14.325 2.87 14.325 2.3 12.2 2.3  ;
        POLYGON 9.295 1.82 10.555 1.82 10.555 3.15 12.26 3.15 12.26 2.53 13.9 2.53 13.9 3.16 14.785 3.16 14.785 1.26 15.015 1.26 15.015 3.16 15.905 3.16 15.905 2.07 16.245 2.07 16.245 3.39 13.67 3.39 13.67 2.765 12.49 2.765 12.49 3.39 10.325 3.39 10.325 2.05 9.13 2.05 9.13 2.86 8.9 2.86 8.9 1.82 9.065 1.82 9.065 0.99 9.405 0.99 9.405 1.275 9.295 1.275  ;
        POLYGON 15.425 0.8 15.675 0.8 15.675 1.54 16.885 1.54 16.885 2.315 18.29 2.315 18.29 1.46 18.63 1.46 18.63 2.55 16.655 2.55 16.655 1.775 15.675 1.775 15.675 2.87 15.425 2.87  ;
        POLYGON 17.2 0.995 18.965 0.995 18.965 0.575 19.195 0.575 19.195 1.565 20.245 1.565 20.245 1.275 20.515 1.275 20.515 2.085 20.245 2.085 20.245 1.795 19.195 1.795 19.195 3.345 18.965 3.345 18.965 1.23 17.45 1.23 17.45 2.08 17.2 2.08  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_2
