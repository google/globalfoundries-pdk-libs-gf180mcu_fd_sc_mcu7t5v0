# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 30.24 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.3545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 22.49 1.765 23.43 1.765 23.43 2.155 22.49 2.155  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.605 1.21 21.14 1.21 21.14 2.19 20.605 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.785 2.385 28.725 2.385 29.255 2.385 29.255 1.535 25.85 1.535 25.85 0.61 26.435 0.61 26.435 1.205 28.135 1.205 28.135 0.61 28.695 0.61 28.695 1.205 29.54 1.205 29.54 2.655 28.725 2.655 28.085 2.655 28.085 3.38 27.585 3.38 27.585 2.655 26.18 2.655 26.18 3.38 25.785 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.395 3.62 13.01 3.62 13.01 3.445 13.35 3.445 13.35 3.62 16.2 3.62 16.2 3.445 16.56 3.445 16.56 3.62 18.275 3.62 20.465 3.62 20.465 2.915 20.695 2.915 20.695 3.62 22.63 3.62 22.63 2.97 22.97 2.97 22.97 3.62 24.49 3.62 24.765 3.62 24.765 2.53 24.995 2.53 24.995 3.62 26.805 3.62 26.805 3 27.035 3 27.035 3.62 28.725 3.62 28.845 3.62 28.845 3 29.075 3 29.075 3.62 30.24 3.62 30.24 4.22 28.725 4.22 24.49 4.22 18.275 4.22 10.395 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 30.24 -0.3 30.24 0.3 29.765 0.3 29.765 0.925 29.535 0.925 29.535 0.3 27.525 0.3 27.525 0.925 27.295 0.925 27.295 0.3 25.285 0.3 25.285 0.925 25.055 0.925 25.055 0.3 22.2 0.3 22.2 1.075 21.86 1.075 21.86 0.3 14.14 0.3 14.14 0.915 13.78 0.915 13.78 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.285 6.835 1.285 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.385 9.835 2.385 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.395 1.8 10.395 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 11.68 2.525 14.6 2.525 14.6 2.78 14.16 2.78 14.16 2.755 12.2 2.755 12.2 2.775 11.68 2.775  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 15.905 2.065 15.905 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 14.96 2.525 16.325 2.525 16.325 1.835 12.295 1.835 12.295 1.605 16.325 1.605 16.325 0.99 16.665 0.99 16.665 2.525 17.79 2.525 17.79 2.78 17.36 2.78 17.36 2.755 15.4 2.755 15.4 2.78 14.96 2.78  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.81 2.985 13.81 3.16 15.74 3.16 15.74 2.985 17.02 2.985 17.02 3.16 18.045 3.16 18.045 2.035 18.275 2.035 18.275 3.39 16.79 3.39 16.79 3.215 15.97 3.215 15.97 3.39 13.58 3.39 13.58 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.37 1.145 14.37 0.53 19.675 0.53 19.675 1.765 19.445 1.765 19.445 0.76 17.17 0.76 17.17 1.745 16.94 1.745 16.94 0.76 14.6 0.76 14.6 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 18.57 0.99 19.215 0.99 19.215 1.995 19.955 1.995 19.955 0.715 21.63 0.715 21.63 1.925 21.77 1.925 21.77 2.93 21.43 2.93 21.43 2.155 21.4 2.155 21.4 0.96 20.185 0.96 20.185 2.225 19.775 2.225 19.775 2.835 19.545 2.835 19.545 2.225 18.985 2.225 18.985 1.22 18.57 1.22  ;
        POLYGON 17.445 0.99 17.785 0.99 17.785 1.575 18.755 1.575 18.755 3.16 20.005 3.16 20.005 2.455 21.155 2.455 21.155 3.16 22.08 3.16 22.08 2.51 23.43 2.51 23.43 3.16 24.26 3.16 24.26 1.91 24.49 1.91 24.49 3.39 23.2 3.39 23.2 2.74 22.315 2.74 22.315 3.39 20.925 3.39 20.925 2.685 20.235 2.685 20.235 3.39 18.525 3.39 18.525 1.805 17.445 1.805  ;
        POLYGON 22.01 1.305 24.335 1.305 24.335 0.655 24.565 0.655 24.565 1.305 25.175 1.305 25.175 1.825 28.725 1.825 28.725 2.095 24.945 2.095 24.945 1.535 24.03 1.535 24.03 2.93 23.69 2.93 23.69 1.535 22.24 1.535 22.24 2.2 22.01 2.2  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
