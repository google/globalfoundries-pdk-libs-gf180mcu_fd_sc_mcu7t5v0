# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.84 1.23 7.18 1.23 7.18 2.33 7.72 2.33 7.72 2.71 6.84 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.14 2.33 5.72 2.33 5.72 1.535 6.04 1.535 6.04 2.71 5.14 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.35 1.77 3.8 1.77 3.8 2.15 2.35 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.04 1.105 4.36 1.105 4.36 1.77 4.95 1.77 4.95 2.15 4.04 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.8 0.55 2.12 0.55 2.12 2.235 1.8 2.235  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.48 1.77 1.24 1.77 1.24 0.55 1.56 0.55 1.56 2.15 0.48 2.15  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7565 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.51 0.55 4.895 0.55 4.895 0.865 5.88 0.865 5.88 0.67 7.635 0.67 7.635 1 6.6 1 6.6 2.77 6.28 2.77 6.28 1.095 4.665 1.095 4.665 0.78 2.51 0.78  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.685 2.53 0.685 3.62 2.44 3.62 2.44 3.04 2.67 3.04 2.67 3.62 7.635 3.62 7.84 3.62 7.84 4.22 7.635 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 5.485 0.3 5.485 0.635 5.145 0.635 5.145 0.3 0.71 0.3 0.71 0.905 0.48 0.905 0.48 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 2.53 4.5 2.53 4.5 2.76 1.705 2.76 1.705 3.38 1.365 3.38  ;
        POLYGON 3.095 3.095 7.635 3.095 7.635 3.325 3.095 3.325  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_1
