# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.612 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.66 5.7 1.66 5.7 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.0968 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.085 2.33 12.805 2.33 13.32 2.33 13.32 1.42 8.085 1.42 8.085 0.675 8.345 0.675 8.345 0.98 10.325 0.98 10.325 0.675 10.555 0.675 10.555 0.98 12.565 0.98 12.565 0.675 12.795 0.675 12.795 0.98 14.805 0.98 14.805 0.675 15.035 0.675 15.035 0.98 17.045 0.98 17.045 0.675 17.275 0.675 17.275 0.98 19.285 0.98 19.285 0.53 19.515 0.53 19.515 1.42 14.12 1.42 14.12 2.33 19.415 2.33 19.415 3.38 19.185 3.38 19.185 2.93 17.175 2.93 17.175 3.38 16.945 3.38 16.945 2.93 14.935 2.93 14.935 3.38 14.705 3.38 14.705 2.93 12.805 2.93 12.695 2.93 12.695 3.38 12.465 3.38 12.465 2.93 10.455 2.93 10.455 3.38 10.225 3.38 10.225 2.93 8.315 2.93 8.315 3.38 8.085 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 2.53 7.095 2.53 7.095 3.62 9.105 3.62 9.105 3.17 9.335 3.17 9.335 3.62 11.345 3.62 11.345 3.17 11.575 3.17 11.575 3.62 12.805 3.62 13.585 3.62 13.585 3.17 13.815 3.17 13.815 3.62 15.825 3.62 15.825 3.17 16.055 3.17 16.055 3.62 18.065 3.62 18.065 3.17 18.295 3.17 18.295 3.62 20.26 3.62 20.305 3.62 20.305 2.53 20.535 2.53 20.535 3.62 21.28 3.62 21.28 4.22 20.26 4.22 12.805 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.69 0.3 20.69 0.765 20.35 0.765 20.35 0.3 18.45 0.3 18.45 0.71 18.11 0.71 18.11 0.3 16.21 0.3 16.21 0.71 15.87 0.71 15.87 0.3 13.97 0.3 13.97 0.71 13.63 0.71 13.63 0.3 11.73 0.3 11.73 0.71 11.39 0.71 11.39 0.3 9.49 0.3 9.49 0.71 9.15 0.71 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 6.26 2.53 6.26 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 5.845 1.015 5.845 0.675 6.075 0.675 6.075 1.015 6.495 1.015 6.495 1.685 12.805 1.685 12.805 2.025 6.495 2.025 6.495 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 14.625 1.685 20.26 1.685 20.26 2.03 14.625 2.03  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_12
