# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 34.72 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 11.02 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.74 9.9 1.74 9.9 2.15 0.63 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.565 2.27 21.57 2.27 22.23 2.27 22.23 1.51 12.565 1.51 12.565 0.675 12.825 0.675 12.825 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 0.865 19.285 0.865 19.285 0.675 19.515 0.675 19.515 0.865 21.525 0.865 21.525 0.675 21.755 0.675 21.755 0.865 23.765 0.865 23.765 0.675 23.995 0.675 23.995 0.865 26.005 0.865 26.005 0.675 26.235 0.675 26.235 0.865 28.245 0.865 28.245 0.675 28.475 0.675 28.475 0.865 30.485 0.865 30.485 0.675 30.715 0.675 30.715 0.865 32.725 0.865 32.725 0.675 32.955 0.675 32.955 1.51 23.13 1.51 23.13 2.27 32.855 2.27 32.855 3.38 32.625 3.38 32.625 3 30.615 3 30.615 3.38 30.385 3.38 30.385 3 28.375 3 28.375 3.38 28.145 3.38 28.145 3 26.135 3 26.135 3.38 25.905 3.38 25.905 3 23.895 3 23.895 3.38 23.665 3.38 23.665 3 21.655 3 21.655 3.38 21.57 3.38 21.425 3.38 21.425 3 19.415 3 19.415 3.38 19.185 3.38 19.185 3 17.175 3 17.175 3.38 16.945 3.38 16.945 3 14.935 3 14.935 3.38 14.705 3.38 14.705 3 12.795 3 12.795 3.38 12.565 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 3 7.095 3 7.095 3.62 9.105 3.62 9.105 3 9.335 3 9.335 3.62 11.345 3.62 11.345 2.53 11.575 2.53 11.575 3.62 13.585 3.62 13.585 3.23 13.815 3.23 13.815 3.62 15.825 3.62 15.825 3.23 16.055 3.23 16.055 3.62 18.065 3.62 18.065 3.23 18.295 3.23 18.295 3.62 20.305 3.62 20.305 3.23 20.535 3.23 20.535 3.62 21.57 3.62 22.545 3.62 22.545 3.23 22.775 3.23 22.775 3.62 24.785 3.62 24.785 3.23 25.015 3.23 25.015 3.62 27.025 3.62 27.025 3.23 27.255 3.23 27.255 3.62 29.265 3.62 29.265 3.23 29.495 3.23 29.495 3.62 31.505 3.62 31.505 3.23 31.735 3.23 31.735 3.62 33.6 3.62 33.745 3.62 33.745 2.53 33.975 2.53 33.975 3.62 34.72 3.62 34.72 4.22 33.6 4.22 21.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 34.72 -0.3 34.72 0.3 34.075 0.3 34.075 1.16 33.845 1.16 33.845 0.3 31.89 0.3 31.89 0.635 31.55 0.635 31.55 0.3 29.65 0.3 29.65 0.635 29.31 0.635 29.31 0.3 27.41 0.3 27.41 0.635 27.07 0.635 27.07 0.3 25.17 0.3 25.17 0.635 24.83 0.635 24.83 0.3 22.93 0.3 22.93 0.635 22.59 0.635 22.59 0.3 20.69 0.3 20.69 0.635 20.35 0.635 20.35 0.3 18.45 0.3 18.45 0.635 18.11 0.635 18.11 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.675 0.3 11.675 0.96 11.445 0.96 11.445 0.3 9.435 0.3 9.435 0.96 9.205 0.96 9.205 0.3 7.195 0.3 7.195 0.96 6.965 0.96 6.965 0.3 4.955 0.3 4.955 0.96 4.725 0.96 4.725 0.3 2.715 0.3 2.715 0.96 2.485 0.96 2.485 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 10.225 2.53 10.225 1.42 1.365 1.42 1.365 0.675 1.595 0.675 1.595 1.19 3.605 1.19 3.605 0.675 3.835 0.675 3.835 1.19 5.845 1.19 5.845 0.675 6.075 0.675 6.075 1.19 8.085 1.19 8.085 0.675 8.315 0.675 8.315 1.19 10.325 1.19 10.325 0.675 10.68 0.675 10.68 1.74 21.57 1.74 21.57 1.97 10.68 1.97 10.68 3.38 10.225 3.38 10.225 2.76 8.215 2.76 8.215 3.38 7.985 3.38 7.985 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.595 2.76 1.595 3.38 1.365 3.38  ;
        POLYGON 23.68 1.74 33.6 1.74 33.6 1.97 23.68 1.97  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_20
