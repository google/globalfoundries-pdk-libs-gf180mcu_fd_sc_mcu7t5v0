* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS
