# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 26.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.62 1.17 20.11 1.17 20.11 2.19 19.62 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0791 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.555 2.38 25.3 2.38 25.53 2.38 25.53 1.535 24.17 1.535 24.17 0.61 24.695 0.61 24.695 1.265 25.795 1.265 25.795 2.655 25.3 2.655 25.1 2.655 25.1 3.38 24.555 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.39 3.62 13.19 3.62 13.19 3.445 13.53 3.445 13.53 3.62 15.46 3.62 15.46 2.91 15.82 2.91 15.82 3.62 17.25 3.62 19.485 3.62 19.485 2.965 19.825 2.965 19.825 3.62 21.58 3.62 21.58 2.965 21.92 2.965 21.92 3.62 22.54 3.62 23.54 3.62 23.54 2.53 23.77 2.53 23.77 3.62 25.3 3.62 25.595 3.62 25.595 2.945 25.825 2.945 25.825 3.62 26.32 3.62 26.32 4.22 25.3 4.22 22.54 4.22 17.25 4.22 10.39 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 26.32 -0.3 26.32 0.3 25.825 0.3 25.825 0.905 25.595 0.905 25.595 0.3 23.545 0.3 23.545 0.905 23.315 0.905 23.315 0.3 21.705 0.3 21.705 0.89 21.475 0.89 21.475 0.3 13.48 0.3 13.48 0.915 13.12 0.915 13.12 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.74 4.63 1.74 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.485 9.835 2.485 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.39 1.8 10.39 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 14.255 2.065 14.255 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 12.475 1.605 14.715 1.605 14.715 1.99 15.47 1.99 15.47 0.99 15.81 0.99 15.81 1.99 16.74 1.99 16.74 2.885 16.51 2.885 16.51 2.22 14.715 2.22 14.715 2.93 14.485 2.93 14.485 1.835 12.475 1.835  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.99 2.985 13.99 3.16 15 3.16 15 2.45 16.28 2.45 16.28 3.115 17.02 3.115 17.02 2.065 17.25 2.065 17.25 3.345 16.05 3.345 16.05 2.68 15.23 2.68 15.23 3.39 13.76 3.39 13.76 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.1 1.145 14.1 0.53 18.82 0.53 18.82 1.815 18.45 1.815 18.45 0.76 16.32 0.76 16.32 1.74 16.09 1.74 16.09 0.76 14.33 0.76 14.33 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 17.71 0.99 18.22 0.99 18.22 2.045 19.05 2.045 19.05 0.53 20.865 0.53 20.865 2.93 20.525 2.93 20.525 0.76 19.28 0.76 19.28 2.275 18.78 2.275 18.78 2.885 18.55 2.885 18.55 2.315 17.99 2.315 17.99 1.265 17.71 1.265  ;
        POLYGON 16.59 0.99 16.93 0.99 16.93 1.525 17.76 1.525 17.76 3.115 19.01 3.115 19.01 2.505 20.285 2.505 20.285 3.16 21.1 3.16 21.1 2.505 22.2 2.505 22.2 1.96 22.54 1.96 22.54 2.735 21.33 2.735 21.33 3.39 20.055 3.39 20.055 2.735 19.24 2.735 19.24 3.345 17.53 3.345 17.53 1.76 16.59 1.76  ;
        POLYGON 21.115 1.495 22.595 1.495 22.595 0.655 23.03 0.655 23.03 1.825 25.3 1.825 25.3 2.095 23.03 2.095 23.03 3.38 22.8 3.38 22.8 1.725 21.345 1.725 21.345 2.17 21.115 2.17  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
