# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.89 1.77 3.895 1.77 3.895 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.3955 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.65 0.65 15.14 0.65 15.14 1.59 14.65 1.59  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 1.575 1.77 1.575 2.15 0.71 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.08 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.38 2.33 20.28 2.33 20.81 2.33 20.81 1.175 18.435 1.175 18.435 0.79 18.665 0.79 18.665 0.945 20.635 0.945 20.635 0.79 21.19 0.79 21.19 2.765 20.76 2.765 20.76 3.235 20.42 3.235 20.42 2.765 20.28 2.765 18.72 2.765 18.72 3.235 18.38 3.235  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.035 3.62 3.17 3.62 3.17 2.845 3.51 2.845 3.51 3.62 5.015 3.62 7.59 3.62 7.59 3.005 7.93 3.005 7.93 3.62 9.17 3.62 9.605 3.62 9.605 2.79 9.835 2.79 9.835 3.62 10.33 3.62 10.855 3.62 14.22 3.62 14.22 3.28 14.56 3.28 14.56 3.62 16.385 3.62 16.595 3.62 16.595 2.69 16.825 2.69 16.825 3.62 17.415 3.62 17.415 2.69 17.645 2.69 17.645 3.62 19.455 3.62 19.455 3.16 19.685 3.16 19.685 3.62 20.28 3.62 21.495 3.62 21.495 2.69 21.725 2.69 21.725 3.62 22.4 3.62 22.4 4.22 20.28 4.22 16.385 4.22 10.855 4.22 10.33 4.22 9.17 4.22 5.015 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.025 0.3 22.025 0.765 21.795 0.765 21.795 0.3 19.84 0.3 19.84 0.715 19.5 0.715 19.5 0.3 17.545 0.3 17.545 0.765 17.315 0.765 17.315 0.3 14.405 0.3 14.405 1.13 14.175 1.13 14.175 0.3 8.87 0.3 8.87 0.915 8.53 0.915 8.53 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 0.915 1.31 0.915 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.465 1.805 2.465 1.805 1.375 0.245 1.375 0.245 0.63 0.475 0.63 0.475 1.145 2.035 1.145 2.035 2.7 0.575 2.7 0.575 2.805 0.345 2.805  ;
        POLYGON 4.245 0.79 4.555 0.79 4.555 2.8 4.245 2.8  ;
        POLYGON 2.615 2.38 4.015 2.38 4.015 3.16 4.785 3.16 4.785 1.555 5.015 1.555 5.015 3.39 3.785 3.39 3.785 2.61 2.615 2.61 2.615 2.805 2.385 2.805 2.385 0.63 2.715 0.63 2.715 0.97 2.615 0.97  ;
        POLYGON 6.285 2.545 8.39 2.545 8.39 2.83 9.17 2.83 9.17 3.06 8.16 3.06 8.16 2.775 6.515 2.775 6.515 3.115 6.285 3.115  ;
        POLYGON 5.265 0.79 5.675 0.79 5.675 2.085 8.85 2.085 8.85 2.24 10.33 2.24 10.33 2.47 8.62 2.47 8.62 2.315 5.495 2.315 5.495 2.8 5.265 2.8  ;
        POLYGON 6.93 1.625 10.09 1.625 10.09 0.99 10.43 0.99 10.43 1.78 10.855 1.78 10.855 3.13 10.625 3.13 10.625 2.01 10.06 2.01 10.06 1.855 6.93 1.855  ;
        POLYGON 6.17 1.165 9.1 1.165 9.1 0.53 12.625 0.53 12.625 2.525 12.395 2.525 12.395 0.76 11.255 0.76 11.255 1.62 11.025 1.62 11.025 0.76 9.33 0.76 9.33 1.395 6.515 1.395 6.515 1.565 6.17 1.565  ;
        POLYGON 12.98 0.82 13.32 0.82 13.32 2.93 12.98 2.93  ;
        POLYGON 11.645 0.99 11.995 0.99 11.995 2.065 12.105 2.065 12.105 3.16 13.67 3.16 13.67 2.815 15.02 2.815 15.02 3.155 16.135 3.155 16.135 2.035 16.385 2.035 16.385 2.375 16.365 2.375 16.365 3.39 14.79 3.39 14.79 3.05 13.9 3.05 13.9 3.39 11.875 3.39 11.875 2.405 11.645 2.405  ;
        POLYGON 13.56 1.77 13.9 1.77 13.9 2.235 15.56 2.235 15.56 1.435 16.595 1.435 16.595 0.74 16.825 0.74 16.825 1.435 20.28 1.435 20.28 1.665 15.79 1.665 15.79 2.87 15.45 2.87 15.45 2.47 13.56 2.47  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
