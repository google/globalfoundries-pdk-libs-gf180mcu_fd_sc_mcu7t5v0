# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.91 1.325 3.495 1.325 3.495 1.17 3.785 1.17 3.785 1.325 5.735 1.325 5.735 1.17 6.105 1.17 6.105 1.59 2.91 1.59  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.53 1.82 5.55 1.82 5.55 2.105 1.53 2.105  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 1.82 1.16 1.82 1.16 2.38 5.945 2.38 5.945 1.82 6.57 1.82 6.57 2.115 6.175 2.115 6.175 2.655 0.87 2.655  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2436 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.315 2.36 11.095 2.36 11.345 2.36 11.345 1.535 8.265 1.535 8.265 0.53 8.495 0.53 8.495 1.265 10.505 1.265 10.505 0.53 10.735 0.53 10.735 1.265 11.62 1.265 11.62 2.68 11.095 2.68 10.685 2.68 10.685 3.39 10.455 3.39 10.455 2.68 8.545 2.68 8.545 3.39 8.315 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 6.865 3.62 6.865 3.06 7.095 3.06 7.095 3.62 9.335 3.62 9.335 3 9.565 3 9.565 3.62 11.095 3.62 11.525 3.62 11.525 3 11.755 3 11.755 3.62 12.32 3.62 12.32 4.22 11.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.855 0.3 11.855 0.97 11.625 0.97 11.625 0.3 9.615 0.3 9.615 0.9 9.385 0.9 9.385 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.005 0.245 1.005 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 3.505 2.935 6.405 2.935 6.405 2.52 6.8 2.52 6.8 1.095 6.36 1.095 6.36 0.92 5.495 0.92 5.495 1.095 4.19 1.095 4.19 0.92 3.26 0.92 3.26 1.095 1.94 1.095 1.94 0.775 1.265 0.775 1.265 0.545 2.185 0.545 2.185 0.865 3.015 0.865 3.015 0.545 4.43 0.545 4.43 0.865 5.26 0.865 5.26 0.545 6.62 0.545 6.62 0.865 7.03 0.865 7.03 1.765 11.095 1.765 11.095 1.995 7.03 1.995 7.03 2.755 6.635 2.755 6.635 3.22 3.505 3.22  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_4
