* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
M_n_tran_1 VSS A ZN VPW nmos_5p0 W=8.2e-07 L=6e-07
M_transistor_0 VDD A A VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
