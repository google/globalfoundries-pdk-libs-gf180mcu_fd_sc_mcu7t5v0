* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latsnq_1 D E SETN Q VDD VNW VPW VSS
M_tn2 net6 E VSS VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn7 VSS D net2 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn6 net3 E net2 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn5 net4 net6 net3 VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn4 net4 net1 VSS VPW nmos_5p0 W=3.95e-07 L=6e-07
M_tn9 VSS net3 net0 VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn8 net0 SETN net1 VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn3 net5 net1 VSS VPW nmos_5p0 W=4.65e-07 L=6e-07
M_tn0 Q net5 VSS VPW nmos_5p0 W=8.2e-07 L=6e-07
M_tp2 net6 E VDD VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp6 VDD D net7 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp5 net7 net6 net3 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp4 net3 E net8 VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp3 net8 net1 VDD VNW pmos_5p0 W=6.3e-07 L=5e-07
M_tp9 VDD net3 net1 VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp8 net1 SETN VDD VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp7 net5 net1 VDD VNW pmos_5p0 W=9.25e-07 L=5e-07
M_tp0 Q net5 VDD VNW pmos_5p0 W=1.22e-06 L=5e-07
.ENDS
