# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.595 1.8 3.5 1.8 3.5 2.12 1.595 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.765 1.21 1.765 1.21 2.36 3.93 2.36 3.93 1.825 4.275 1.825 4.275 2.68 0.87 2.68  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.085 2.36 8.96 2.36 9.205 2.36 9.205 1.54 5.985 1.54 5.985 0.53 6.215 0.53 6.215 1.26 8.225 1.26 8.225 0.53 8.455 0.53 8.455 1.265 9.46 1.265 9.46 2.68 8.96 2.68 8.405 2.68 8.405 3.39 8.175 3.39 8.175 2.68 6.315 2.68 6.315 3.39 6.085 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.965 3.62 4.965 2.53 5.195 2.53 5.195 3.62 7.105 3.62 7.105 2.935 7.335 2.935 7.335 3.62 8.96 3.62 9.245 3.62 9.245 2.94 9.475 2.94 9.475 3.62 10.08 3.62 10.08 4.22 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.575 0.3 9.575 0.98 9.345 0.98 9.345 0.3 7.335 0.3 7.335 0.985 7.105 0.985 7.105 0.3 4.955 0.3 4.955 1.07 4.725 1.07 4.725 0.3 2.715 0.3 2.715 1.07 2.485 1.07 2.485 0.3 0.475 0.3 0.475 1.07 0.245 1.07 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.35 2.945 4.505 2.945 4.505 1.57 1.365 1.57 1.365 0.53 1.595 0.53 1.595 1.325 3.605 1.325 3.605 0.53 3.835 0.53 3.835 1.325 4.735 1.325 4.735 1.825 8.96 1.825 8.96 2.095 4.735 2.095 4.735 3.215 2.35 3.215  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_4
