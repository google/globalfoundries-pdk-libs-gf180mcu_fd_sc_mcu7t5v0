# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.58 1.8 18.44 1.8 18.44 2.12 14.58 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.29 1.76 19.53 1.76 19.53 2.36 22.6 2.36 22.6 1.92 23.96 1.92 23.96 2.36 27.25 2.36 27.25 1.76 27.49 1.76 27.49 2.59 24.605 2.59 24.605 2.71 21.955 2.71 21.955 2.59 19.29 2.59  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.18 1.8 21.685 1.8 21.685 1.45 24.775 1.45 24.775 1.8 26.835 1.8 26.835 2.12 24.545 2.12 24.545 1.68 21.915 1.68 21.915 2.12 20.18 2.12  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.58 1.8 13.34 1.8 13.34 2.12 9.58 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.775 1.53 1.095 1.53 1.095 2.36 4.16 2.36 4.16 1.92 5.52 1.92 5.52 2.36 8.58 2.36 8.58 1.76 8.84 1.76 8.84 2.595 6.16 2.595 6.16 2.7 3.52 2.7 3.52 2.595 0.775 2.595  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.74 1.8 3.59 1.8 3.59 1.335 6.45 1.335 6.45 1.8 8.31 1.8 8.31 2.12 6.22 2.12 6.22 1.565 3.82 1.565 3.82 2.12 1.74 2.12  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.0289 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.58 2.36 13.57 2.36 13.57 0.99 26.82 0.99 26.82 1.22 13.87 1.22 13.87 2.36 17.89 2.36 17.89 2.795 9.58 2.795  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.285 2.77 3.285 2.77 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 13.87 3.62 20.87 3.62 20.87 3.285 21.21 3.285 21.21 3.62 25.35 3.62 25.35 3.285 25.69 3.285 25.69 3.62 27.995 3.62 28.16 3.62 28.56 3.62 28.56 4.22 28.16 4.22 27.995 4.22 13.87 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 28.56 -0.3 28.56 0.3 12.85 0.3 12.85 0.635 12.51 0.635 12.51 0.3 10.61 0.3 10.61 0.635 10.27 0.635 10.27 0.3 8.37 0.3 8.37 0.635 8.03 0.635 8.03 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.295 2.53 0.525 2.53 0.525 2.825 3.27 2.825 3.27 3.09 6.41 3.09 6.41 2.825 7.73 2.825 7.73 3.09 13.87 3.09 13.87 3.32 7.5 3.32 7.5 3.055 6.66 3.055 6.66 3.32 3.02 3.32 3.02 3.055 0.525 3.055 0.525 3.38 0.295 3.38  ;
        POLYGON 14.24 3.09 20.11 3.09 20.11 2.825 21.705 2.825 21.705 3.09 24.855 3.09 24.855 2.825 27.765 2.825 27.765 2.53 27.995 2.53 27.995 3.38 27.765 3.38 27.765 3.055 25.1 3.055 25.1 3.32 21.46 3.32 21.46 3.055 20.355 3.055 20.355 3.32 14.24 3.32  ;
        POLYGON 0.18 0.865 13.1 0.865 13.1 0.53 28.16 0.53 28.16 0.76 13.33 0.76 13.33 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_4
