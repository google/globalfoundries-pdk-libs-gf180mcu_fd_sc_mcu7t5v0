# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.62 1.1 1.06 1.1 1.06 1.715 2.15 1.715 2.15 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3656 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.605 2.36 4.095 2.36 4.36 2.36 4.36 1.42 3.605 1.42 3.605 0.675 3.865 0.675 3.865 1.14 5.845 1.14 5.845 0.675 6.075 0.675 6.075 1.42 5.16 1.42 5.16 2.36 5.975 2.36 5.975 3.38 5.745 3.38 5.745 2.68 4.095 2.68 3.835 2.68 3.835 3.38 3.605 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.095 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.81 3.62 6.865 3.62 6.865 2.57 7.095 2.57 7.095 3.62 7.84 3.62 7.84 4.22 6.81 4.22 4.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 2.53 2.67 2.53 2.67 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 2.905 1.015 2.905 1.685 4.095 1.685 4.095 2.025 2.905 2.025 2.905 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 5.585 1.685 6.81 1.685 6.81 2.025 5.585 2.025  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_4
