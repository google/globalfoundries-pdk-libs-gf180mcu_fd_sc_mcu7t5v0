# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.05 1.77 4.05 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.38 1.77 20.63 1.77 20.63 2.15 19.38 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1495 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 18.225 1.77 18.225 1.34 18.54 1.34 18.54 2.15 17.45 2.15  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.15 0.28 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0582 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.545 2.07 23.72 2.07 24.17 2.07 24.17 1.17 23.6 1.17 23.6 0.55 23.98 0.55 23.98 0.94 24.55 0.94 24.55 2.32 23.98 2.32 23.98 3.38 23.72 3.38 23.545 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.055 3.62 3.05 3.62 3.05 3 3.39 3 3.39 3.62 7.585 3.62 7.585 3.165 7.93 3.165 7.93 3.62 13.45 3.62 13.45 3.035 13.68 3.035 13.68 3.62 15.48 3.62 17.705 3.62 17.705 2.94 18.045 2.94 18.045 3.62 19.745 3.62 19.745 2.94 20.085 2.94 20.085 3.62 21.61 3.62 21.84 3.62 21.84 2.415 22.07 2.415 22.07 3.62 22.58 3.62 22.58 2.57 22.81 2.57 22.81 3.62 23.72 3.62 24.62 3.62 24.62 2.57 24.85 2.57 24.85 3.62 25.2 3.62 25.2 4.22 23.72 4.22 21.61 4.22 15.48 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 25.005 0.3 25.005 0.71 24.665 0.71 24.665 0.3 22.71 0.3 22.71 0.765 22.48 0.765 22.48 0.3 20.085 0.3 20.085 1.075 19.745 1.075 19.745 0.3 10.92 0.3 10.92 0.915 10.58 0.915 10.58 0.3 3.61 0.3 3.61 1.075 3.27 1.075 3.27 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.435 1.825 2.435 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.67 0.575 2.67 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 0.845 4.73 0.845 4.73 2.83 4.29 2.83  ;
        POLYGON 6.405 2.245 8.97 2.245 8.97 2.585 10.85 2.585 10.85 2.875 10.51 2.875 10.51 2.815 8.74 2.815 8.74 2.475 6.635 2.475 6.635 2.87 6.405 2.87  ;
        POLYGON 5.31 1.785 5.565 1.785 5.565 0.79 5.795 0.79 5.795 1.785 9.43 1.785 9.43 2.07 12.07 2.07 12.07 1.545 12.47 1.545 12.47 1.775 12.3 1.775 12.3 2.3 9.2 2.3 9.2 2.015 5.65 2.015 5.65 2.83 5.31 2.83  ;
        POLYGON 11.79 2.645 12.53 2.645 12.53 2.115 14.465 2.115 14.465 1.315 11.84 1.315 11.84 1.835 9.66 1.835 9.66 1.555 7.03 1.555 7.03 1.325 9.89 1.325 9.89 1.605 11.61 1.605 11.61 1.085 14.75 1.085 14.75 2.125 14.975 2.125 14.975 2.875 14.635 2.875 14.635 2.345 12.76 2.345 12.76 2.875 11.79 2.875  ;
        POLYGON 2.615 2.54 4.015 2.54 4.015 3.105 6.865 3.105 6.865 2.705 8.51 2.705 8.51 3.16 12.99 3.16 12.99 2.575 14.405 2.575 14.405 3.16 15.25 3.16 15.25 2.07 15.48 2.07 15.48 3.39 14.175 3.39 14.175 2.805 13.22 2.805 13.22 3.39 8.28 3.39 8.28 2.935 7.095 2.935 7.095 3.335 3.785 3.335 3.785 2.77 2.615 2.77 2.615 3.3 2.385 3.3 2.385 0.81 2.715 0.81 2.715 1.15 2.615 1.15  ;
        POLYGON 6.135 0.79 10.35 0.79 10.35 1.145 11.15 1.145 11.15 0.53 17.115 0.53 17.115 0.855 16.775 0.855 16.775 0.76 14.77 0.76 14.77 0.855 14.43 0.855 14.43 0.76 11.38 0.76 11.38 1.375 10.12 1.375 10.12 1.02 6.475 1.02 6.475 1.555 6.135 1.555  ;
        POLYGON 16.17 1.03 16.455 1.03 16.455 1.085 17.71 1.085 17.71 0.79 19.01 0.79 19.01 2.855 18.78 2.855 18.78 1.075 17.995 1.075 17.995 1.315 17.015 1.315 17.015 2.895 16.675 2.895 16.675 1.37 16.17 1.37  ;
        POLYGON 14.98 1.085 15.94 1.085 15.94 3.16 17.245 3.16 17.245 2.475 18.505 2.475 18.505 3.085 19.24 3.085 19.24 2.48 20.545 2.48 20.545 3.085 21.38 3.085 21.38 1.91 21.61 1.91 21.61 3.32 20.315 3.32 20.315 2.71 19.47 2.71 19.47 3.32 18.275 3.32 18.275 2.71 17.475 2.71 17.475 3.39 15.71 3.39 15.71 1.315 14.98 1.315  ;
        POLYGON 20.82 2.515 20.92 2.515 20.92 1.54 19.305 1.54 19.305 1.31 21.76 1.31 21.76 0.79 21.99 0.79 21.99 1.33 23.305 1.33 23.305 1.475 23.72 1.475 23.72 1.82 22.965 1.82 22.965 1.56 21.15 1.56 21.15 2.855 20.82 2.855  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
