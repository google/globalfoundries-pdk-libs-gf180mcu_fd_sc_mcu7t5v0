# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5235 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.77 6.07 1.77 6.07 2.12 4.01 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5235 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.33 1.21 2.71 1.21 2.71 2.71 2.33 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.047 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 1.445 3.295 1.445 3.295 2.36 6.09 2.36 6.09 2.785 2.94 2.785  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 0.65 0.575 0.65 0.575 3.27 0.13 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 2.76 1.595 2.76 1.595 3.62 3.89 3.62 5.31 3.62 5.31 3.105 5.65 3.105 5.65 3.62 6.815 3.62 7.28 3.62 7.28 4.22 6.815 4.22 3.89 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 5.695 0.3 5.695 0.88 5.465 0.88 5.465 0.3 1.595 0.3 1.595 0.865 1.365 0.865 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.055 3.11 3.89 3.11 3.89 3.34 1.825 3.34 1.825 1.625 0.84 1.625 0.84 1.39 1.825 1.39 1.825 0.575 3.88 0.575 3.88 0.815 2.055 0.815  ;
        POLYGON 4.125 1.145 6.35 1.145 6.35 0.53 6.815 0.53 6.815 3.38 6.35 3.38 6.35 1.375 4.125 1.375  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_1
