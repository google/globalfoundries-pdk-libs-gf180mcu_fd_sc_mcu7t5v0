# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.726 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.55 1.08 0.55 1.08 1.74 1.65 1.74 1.65 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0086 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.665 2.36 3.21 2.36 3.47 2.36 3.47 1.51 2.665 1.51 2.665 0.8 2.895 0.8 2.895 1.28 3.81 1.28 3.81 2.71 3.21 2.71 2.895 2.71 2.895 3.39 2.665 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.36 3.62 1.36 3.05 1.7 3.05 1.7 3.62 3.21 3.62 3.685 3.62 3.685 3.05 3.915 3.05 3.915 3.62 4.48 3.62 4.48 4.22 3.21 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 4.07 0.3 4.07 1.05 3.73 1.05 3.73 0.3 1.83 0.3 1.83 1.095 1.49 1.095 1.49 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.805 0.475 0.805 0.475 2.59 1.89 2.59 1.89 1.74 3.21 1.74 3.21 2.04 2.215 2.04 2.215 2.82 0.475 2.82 0.475 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
