# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 1.24 3.31 1.24 3.31 1.56 1.16 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.42 1.8 3.77 1.8 3.77 2.12 0.42 2.12  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.8 5.22 1.8 5.22 2.36 7.885 2.36 7.885 1.8 9.025 1.8 9.025 2.12 8.43 2.12 8.43 2.595 5.665 2.595 5.665 2.71 4.6 2.71  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.65 1.8 7.395 1.8 7.395 2.12 5.65 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1268 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 2.36 4.04 2.36 4.04 1.56 3.655 1.56 3.655 1 2.15 1 2.15 0.68 3.915 0.68 3.915 1.24 4.915 1.24 4.915 0.87 5.41 0.87 5.41 0.56 5.75 0.56 5.75 0.87 7.65 0.87 7.65 0.56 7.99 0.56 7.99 1.1 5.145 1.1 5.145 1.56 4.36 1.56 4.36 2.78 1.17 2.78  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 6.45 3.62 6.45 3.285 6.79 3.285 6.79 3.62 8.955 3.62 9.52 3.62 9.52 4.22 8.955 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.055 0.3 9.055 0.695 8.825 0.695 8.825 0.3 6.87 0.3 6.87 0.64 6.53 0.64 6.53 0.3 4.395 0.3 4.395 0.69 4.165 0.69 4.165 0.3 0.475 0.3 0.475 0.91 0.245 0.91 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.5 0.475 2.5 0.475 3.16 5.91 3.16 5.91 2.825 8.725 2.825 8.725 2.5 8.955 2.5 8.955 3.39 8.725 3.39 8.725 3.055 6.14 3.055 6.14 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_2
