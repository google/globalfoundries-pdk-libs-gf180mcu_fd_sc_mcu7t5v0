# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.545 1.78 1.63 1.78 1.63 2.265 0.545 2.265  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0795 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.92 1.815 6.085 1.815 6.085 2.235 4.92 2.235  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0374 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.805 0.6 7.16 0.6 7.16 3.38 6.805 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.83 3.62 5.83 3.22 6.17 3.22 6.17 3.62 6.565 3.62 7.87 3.62 7.87 2.53 8.21 2.53 8.21 3.62 8.4 3.62 8.4 4.22 6.565 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 8.155 0.3 8.155 0.9 7.925 0.9 7.925 0.3 5.915 0.3 5.915 0.9 5.685 0.9 5.685 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.42 2.78 1.9 2.78 1.9 1.325 0.19 1.325 0.19 0.865 0.53 0.865 0.53 1.095 2.13 1.095 2.13 2.235 3.65 2.235 3.65 2.52 2.13 2.52 2.13 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 5.355 0.53 5.355 1.355 6.51 1.355 6.51 1.585 5.125 1.585 5.125 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.7 3.16 4.46 3.16 4.46 1.545 3.77 1.545 3.77 0.99 4.11 0.99 4.11 1.315 4.69 1.315 4.69 2.7 6.335 2.7 6.335 1.9 6.565 1.9 6.565 2.93 5.175 2.93 5.175 3.39 2.7 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_2
