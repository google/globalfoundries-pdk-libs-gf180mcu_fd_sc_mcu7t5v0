# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 1.24 4 1.24 4 0.55 4.43 0.55 4.43 1.56 3.35 1.56  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.736 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.8 2.15 1.8 2.15 2.75 1.77 2.75 1.77 2.12 0.825 2.12  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.66 0.53 11.08 0.53 11.08 3.38 10.66 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.05 1.595 3.05 1.595 3.62 2.36 3.62 3.485 3.62 3.485 3.085 3.715 3.085 3.715 3.62 5.1 3.62 7.41 3.62 7.41 2.805 7.75 2.805 7.75 3.62 9.17 3.62 9.705 3.62 9.705 2.53 9.935 2.53 9.935 3.62 11.745 3.62 11.745 2.53 11.975 2.53 11.975 3.62 12.32 3.62 12.32 4.22 9.17 4.22 5.1 4.22 2.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 12.075 0.3 12.075 1.055 11.845 1.055 11.845 0.3 9.835 0.3 9.835 1.055 9.605 1.055 9.605 0.3 7.995 0.3 7.995 0.895 7.765 0.895 7.765 0.3 3.615 0.3 3.615 0.825 3.385 0.825 3.385 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.575 0.53 0.575 1.16 2.36 1.16 2.36 1.39 0.575 1.39 0.575 3.39 0.19 3.39  ;
        POLYGON 3.125 2.335 5.1 2.335 5.1 2.565 3.125 2.565  ;
        POLYGON 2.61 0.53 2.95 0.53 2.95 1.855 4.785 1.855 4.785 1.01 5.015 1.01 5.015 1.855 5.985 1.855 5.985 2.81 5.755 2.81 5.755 2.085 2.895 2.085 2.895 3.39 2.61 3.39  ;
        POLYGON 5.1 3.14 6.275 3.14 6.275 0.76 5.2 0.76 5.2 0.53 6.505 0.53 6.505 1.245 8.58 1.245 8.58 1.475 6.505 1.475 6.505 3.37 5.1 3.37  ;
        POLYGON 6.82 2.075 8.83 2.075 8.83 0.53 9.17 0.53 9.17 2.305 8.715 2.305 8.715 3.225 8.485 3.225 8.485 2.305 6.82 2.305  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_2
