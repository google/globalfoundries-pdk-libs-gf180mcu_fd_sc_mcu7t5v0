# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.76 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.477 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.125 1.77 11.48 1.77 11.48 2.15 5.125 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.2244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.63 2.53 17.49 2.53 17.9 2.53 17.9 1.135 12.73 1.135 12.73 0.865 24.27 0.865 24.27 1.135 18.5 1.135 18.5 2.53 23.17 2.53 23.17 3.38 22.83 3.38 22.83 2.97 21.13 2.97 21.13 3.38 20.79 3.38 20.79 2.97 19.09 2.97 19.09 3.38 18.75 3.38 18.75 2.97 17.49 2.97 17.05 2.97 17.05 3.38 16.71 3.38 16.71 2.97 15.01 2.97 15.01 3.38 14.67 3.38 14.67 2.97 12.97 2.97 12.97 3.38 12.63 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.49 3.62 5.49 3.04 5.83 3.04 5.83 3.62 7.53 3.62 7.53 3.04 7.87 3.04 7.87 3.62 9.57 3.62 9.57 3.04 9.91 3.04 9.91 3.62 11.61 3.62 11.61 3.04 11.95 3.04 11.95 3.62 13.65 3.62 13.65 3.285 13.99 3.285 13.99 3.62 15.69 3.62 15.69 3.285 16.03 3.285 16.03 3.62 17.49 3.62 17.73 3.62 17.73 3.285 18.07 3.285 18.07 3.62 19.77 3.62 19.77 3.285 20.11 3.285 20.11 3.62 21.81 3.62 21.81 3.285 22.15 3.285 22.15 3.62 23.705 3.62 23.85 3.62 23.85 3.04 24.19 3.04 24.19 3.62 25.76 3.62 25.76 4.22 23.705 4.22 17.49 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.76 -0.3 25.76 0.3 25.39 0.3 25.39 0.635 25.05 0.635 25.05 0.3 23.15 0.3 23.15 0.635 22.81 0.635 22.81 0.3 20.91 0.3 20.91 0.635 20.57 0.635 20.57 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.19 0.3 14.19 0.635 13.85 0.635 13.85 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.905 2.78 1.905 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.135 1.095 2.135 2.235 3.65 2.235 3.65 2.52 2.135 2.52 2.135 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 5.945 0.705 5.945 0.865 12.01 0.865 12.01 1.365 16.875 1.365 16.875 1.595 11.78 1.595 11.78 1.095 5.695 1.095 5.695 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.685 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.53 11.78 2.53 11.78 1.965 17.49 1.965 17.49 2.195 12.01 2.195 12.01 2.76 10.93 2.76 10.93 3.38 10.59 3.38 10.59 2.76 8.89 2.76 8.89 3.38 8.55 3.38 8.55 2.76 6.85 2.76 6.85 3.38 6.51 3.38 6.51 2.76 4.825 2.76 4.825 3.39 2.685 3.39  ;
        POLYGON 19.01 1.365 23.705 1.365 23.705 1.595 19.01 1.595  ;
        POLYGON 19.33 1.965 23.705 1.965 23.705 2.195 19.33 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_12
