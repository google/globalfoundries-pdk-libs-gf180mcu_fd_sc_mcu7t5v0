# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.45 1.8 7.175 1.8 7.175 2.13 0.45 2.13  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.24 3.545 1.24 3.545 1.325 5.265 1.325 5.265 1.24 7.635 1.24 7.635 1.825 8.11 1.825 8.11 2.095 7.405 2.095 7.405 1.57 0.61 1.57  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2401 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 8.34 2.36 8.34 1.575 7.885 1.575 7.885 1.01 5.035 1.01 5.035 1.095 3.775 1.095 3.775 1.01 2.14 1.01 2.14 0.68 4.005 0.68 4.005 0.865 4.805 0.865 4.805 0.68 8.115 0.68 8.115 1.345 8.57 1.345 8.57 2.68 7.615 2.68 7.615 3.39 7.385 3.39 7.385 2.68 5.575 2.68 5.575 3.39 5.345 3.39 5.345 2.68 3.535 2.68 3.535 3.39 3.305 3.39 3.305 2.68 1.495 2.68 1.495 3.39 1.265 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.285 3.62 2.285 2.93 2.515 2.93 2.515 3.62 4.325 3.62 4.325 2.93 4.555 2.93 4.555 3.62 6.365 3.62 6.365 2.93 6.595 2.93 6.595 3.62 8.405 3.62 8.405 2.93 8.635 2.93 8.635 3.62 8.96 3.62 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 8.69 0.3 8.69 0.635 8.35 0.635 8.35 0.3 4.575 0.3 4.575 0.635 4.235 0.635 4.235 0.3 0.555 0.3 0.555 0.905 0.325 0.905 0.325 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_4
